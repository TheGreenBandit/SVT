   9��?     �9                              �+�           ?�R@�z�
?+�        ´  