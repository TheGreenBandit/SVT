   9�'T                                      �;�P            ���Ϳ��?�z�              ^�AF-       	    ���                      ��AF-           ���                      �AF-       
    ���                      ��AF-           ���                      ���_�            ����?�Q�>�p�@� 2�  C4    ���_�            >���?�Q�>�p�@� 2�  C4  