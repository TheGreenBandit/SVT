   9��?    �fP                              ?���$                   A~�G              ����$                    @��    �4  A�  