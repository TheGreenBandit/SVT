   ���                                      +}��                    >���            