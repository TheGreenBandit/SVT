   �O�     �                               _=f�M           >u>�>�fa    B�  B�    �=f�M           �k�$>�>�fa    B�  ´    ]=f�M           ��(��<�    ´  ´    �=f�M           <����<�    B�  ´    �=f�M           >Ǯ��<�    B�  Ç    �8�f           ����Y��>�)              �8�f           ����Y��?
D              ��8�f           >��Y��?
D              ��8�f           >��Y��>�G�              	��Dj       	               �4      B�    ��Dj       	   �u        �4      B�    ���Dj       
   �u        �4      B�    #��Dj       
   <�        �4      B�    |��Dj          <�        �4      B�    ���Dj          ��Q�        �4      B�    5��Dj          �&fa        �4      B�    ��Dj          �&fa        �4      B�    9��Dj          �Z        �4      B�    ���Dj          ��        �4      B�    �Ȗ0�           ��?xQ�?h��        B�    Ȗ0�           =�G�?xQ�?h��        B�    ���Dj          ����        �4      B�    x���^              @@              C4    ����^              ����@Q�@�      C4  