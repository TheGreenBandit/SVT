   �As    b                              :H6��           �Y    �\(�        C4  