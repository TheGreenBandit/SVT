   �]�     �                              �]�                           ��        <ȟ�                                     !�]�                           �         �]�                           �p        7�]�                                    �]�                           A�        Y�]�                           B         f�]�                           Bp        ��]�                           B�        c�8�f               �
=p>��               X�8�f               �
=p=u�B              =�8�f           ��  @��L�A�            @�V                �`?u    ô        T7���           ?=p����?}p�    ��33      7���           �:�6���?�fn    ��33      m7���           ���	���$?(��    ��33       7���           ?��ֿ��?�,    ��33    