   �)��    Ca2                              RSy�c           ��=q>B�]��=q              ���^              @               �4  