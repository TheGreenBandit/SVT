   � �^                                      ��oG            �.{�.{��(���      C4    ��oG                �
=m��fb��      C4    ��oG            <���.{��(���      C4    ��oG            �.{��\&��z��      C4    f��X       	    ���	                B�    ���X       
    ���	                B�    ���X           ��8                B�    =��X           �Ǯ                B�  