   q��                                       }��           ���
    >��              �a/�           �#�
                      �a/�                                      �a/�           ����33��              5�V           >L��?�  2�  �� @@  B�33  *2??@           �aG�>L�ξ��        ¯�  >s��                                      >s��          >���?z�H���2    ?�  Ç�