   c"��                                     I|{B           A`      �Y        Cx    \|{B           A`  >8Q�A���        C�    m|{B           A`  >�=qBz�        C��   l|{B           A`  >�p�BJ�        C�  