   �y��    O��                              �3�+��           ���>�=q���@        ´    � 8���            �Ǯ    ��        �4    �Tm�x�            =�G��W
?��fb        ´    ZMm�x�            >�??����fb        ´    �m�x�            �p��??����fb        ´    p_m�x�            �nq�aG���fb        ´    �U7�a            ��(�>Y>k�!              �%�p`,            �J=i>����    �4  ´    �+�p`,            ��>����    �4  Ç    ]m�x�            �u�aG���fb        ´    }m�x�            �}p��aG���fb        ´    �Hm�x�            �xQ�??����fb        ´    Km�x�            ���??����fb        ´    Pdm�x�            >#�
??����fb        ´    jNm�x�            >B�]??����fb        ´    �^m�x�            >\(�W
?��fb        ´    zLm�x�            >.{�W
?��fb        ´    	*�8�f            �끿\%��f`    ��  �4    ,�8�f            �
9?����G�    ��  ô    ��8�f            �u�\%��f`    ��  �4    �q�8�f            ��z�?����G�    ��  ô    1 ���^          �z�@�Q�            �4  