   9��?                                      �9��?                                A�    �9��?                                Bp    	9��?                                B�    �9��?                                B�    �9��?                                C    �9��?                                C4    �9��?                                CR    �9��?                                Cp    49��?                                C�    �9��?                                C�    %	9��?                                C�  