    ���     ?G                              �	��Dj       	                       B�    �	��Dj       	   >�=q                B�    �	��Dj       	   ��=r                C�    X��Dj          ��=r                C�    �	��Dj          �
=l                C�    ���Dj          3�                  C�    K��Dj          >�=t                C�    �	��Dj          ?�                B�    �	Ȗ0�           ���?�  ���<#�
    B�    DȖ0�           ?�?�  ���<#�
    B�    P��E�                �Qhh>�\)�   Ç        �	����            �#�
�(�>���B�      A    �
����            =L�ƿ(�>���B�      ��  