   ��\�                                      �	}��                >.{>8Q�              �	��Dj       	    ����                B�    �	��Dj       
    ����                B�    
��Dj           ����                B�    <	��Dj           ����                B�    (	��Dj           ����                B�    N	��Dj           ����                B�  