   2,��                                      &���                <#��Ƨ�              *%Z_�       	    �L��                C�    +%Z_�       
    �L��                C�    ,%Z_�          ��31                C�    -%Z_�          ��z                C�    /���v           =�G��#�:>u´            0���v           >�=q=���>aG�´            1���v           ?�G��#�>aG�´            2���v           ?�=i=�G�>L��´            3���v           ?���=���\(´            4���v           ?�z�=����´            5���v           >W
D�u��´            6���v           =��ռ���\(´            A����               >.{�#�              C����           ��Q�?\(=qB�      B�    D����           ?�?\(=qB�      C�    E����                @�Ͼ��    B�  B�  