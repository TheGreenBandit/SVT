   ���     �x                              �}��                                      �Ȗ0�           ��>B�]>B�]        B�    �Ȗ0�           ?�3/>B�]>B�`        B�    �Ȗ0�           ?L��?�Q�?
>        B�    �Ȗ0�           �#��?�Q�?
>        B�    ��v'&          @   �0(�@�  ��      ?�    ��v'&          @!G��  A�  �      ?�    ����v           �.u?��V<#��®            ����v           ��?Ǯ�#�:®            ����v           ?�?Ǯ�#�:®            ����v           ?0��?��V<#��®            �7���                ?�Q潸Q��p            ���X       	    ���                B�    ���X       
    ���                B�    ���X           ���                B�    ���X           ���                B�    �@��            >�=q>W
>?�X��  �l        �@��            ��=r>W
>?�X��  �l      