   	�(U    -V3                              �M`|�               �6f]�p��        C4    ��|J               ���c�        �4    �P���               @�                    �P���           ��  @�              B4    |P���           @�  @�              �4    �i�3�           @�  ?�fa�p��        �p    i�3�           ��  ?�fa�p��        Bp    }i�3�           �   @����p��        A�    i�3�           @   @����p��        ��  