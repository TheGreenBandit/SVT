   ���     ]�S                              E}��                                      GȖ0�           ��>B�]>B�]        B�    �Ȗ0�           ?�3/>B�]>B�`        B�    �Ȗ0�           ?L��?�Q�?
>        B�    
Ȗ0�           �#��?�Q�?
>        B�    ~���v           �.u?��V<#��®            ����v           ��?Ǯ�#�:®            p���v           ?�?Ǯ�#�:®            ���v           ?0��?��V<#��®            7���                ?�Q潸Q��p            ���X       	    ���                B�    ���X       
    ���                B�    ���X           ���                B�    ���X           ���                B�    �@��            >�=q>W
>?�X��  �l        V@��            ��=r>W
>?�X��  �l        �7���                �G�<�ز�@            ��y�e                ��_    ´            2�ާ(                    BX  �4      C  