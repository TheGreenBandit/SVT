   9��?    >��                              5�$�                    ?�                s�$�                    ?�          B    |�$�                    ?�          B�    Z�$�                    ?�          B�    H�$�                    ?�          C    i�$�                    ?�          C/    n�$�                    ?�          CR    
�$�                    ?�          Cu    3�$�                    ?�          C�    x�$�                    ?�          C��   M�$�                    ?�      �4  C��   ��$�                    ?�      �4  C�    -�$�                    ?�      �4  Cu    w�$�                    ?�      �4  CR    ��$�                    ?�      �4  C/    ��$�                    ?�      �4  C    ��$�                    ?�      �4  B�    ��$�                    ?�      �4  B�    u�$�                    ?�      �4  B    ��$�                    ?�      �4      