   Pѫ     a��                              �CK�|               �������B        B�  