   �O�     =�                              hpJ               �p��@��              ��c'�           ?@     @��        B�    ��c'�           �G�4(  @��        ��   �pJ               ?\(�@��        C4    n��Dj       	   ��M                ´    ���Dj       
   ��M                ´    ��Dj          ��M                ´    ���Dj          ��M                ´  