   9��?                                     �w��       
    Bo��    C3    C4  C  