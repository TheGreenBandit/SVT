   {~V�                                      <{~V�           ����                      P{~V�            �������?�(�´            ]{~V�            �������@�
>´            \{~V�            �������@�
>´            ^{~V�                ���?�(�´            _{~V�                ���@�
>´            `{~V�                ���@�
>´            a{~V�            �   ���A:�M�4  ¬  ´    b{~V�            �Ffb���A:�M    ¬  ´    c{~V�            �^u���Ax��B�  ¬  ´    d{~V�            ��\.���Ax��B�  ¬  ´    W{~V�            ��\.���A��B�  ¬  ´    R{~V�            �W����A��B�  ¬  ´    f{~V�            ��=k���A��;    ¬  ´    Y{~V�            ��S��Q�A��;    ³����    h{~V�            �J�_?��A��;    ³���.    j{~V�            ?������A��;C4  ´  ´    X{~V�            @ʏZ�\A��;    ³���    p{~V�            @�(�@=p�A��;    B� �.    k����            ��  �Y��A�fg�(            i����            �l���Y��A�fg�(            s����            �  �Y��Aٙ��(          