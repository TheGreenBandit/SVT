   c"��    
�u                              4����                                     5����                       ��            6����                       ��            7����                       �)            8����                       �)      �     9����                       �)      B   