   ��                                      �:��           �^�R                      �8}��           <#��=�\(=�              �?}��           �ff^=L��=�              �=��Dj       
                       Ç    �:��Dj       
   ����                Ç    Y5��Dj          ����                Ç    n4��Dj          ���                Ç    ^5��Dj       	   ���                Ç    �:��Dj       	   �^�X                Ç    �:��Dj          ����                Ç    H6��Dj          ��35                Ç    R<Ȗ0�           >���?�
7=��        B�    	;Ȗ0�           ���A?�
7=��        B�    $>����            ��(�(�?&fa        C4    |<��Dj       	   ��Q�                Ç  