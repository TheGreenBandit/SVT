   Z���     W�                              p�b��           ��35��                    q�b��           ?�����                    rP�!�               �1늾#�        B�    s�b��           ������                    t���           ����?��V        C4    u���           ?�3)�̰?�)        �4    v�            ���@�z����k    ��  ¼    w+�z            @0�ؿ�낾�B�      B�    x+�z            @0�������B�      B�    yҽ��           =L���$zп˅"A�            z+�z            �1G������B�      ´    {+�z            �1G������B�      ´    |ҽ��           ?
9��>R����A�      �4    }ҽ��           �#��L�����A�      �4    ~���^           =�Q�@�������A   �  CE    ���^           >��@�fN����A   B  C    ����^           ?�(�@�fN����A   ��  CC    ����^           �Tz�@�fN��\!A  B  C    �����                ?�?�p�        C4    ��܇           �2�]� �\(�              ��܇           �2�]���\(�              ��܇           @,�����\(�              ��܇           @,���� �\(�            