   q��     <�                              OȖ0�            ���@   >��         B�    RȖ0�            ?�Y@   >��         B�    YȖ0�            ?��>��>�         B�    _Ȗ0�            ���>��>�         B�    P7���               �fg?332        B�    .@��                >��U?0��Cl�4          a@��            >���>��U?0��Cl�4          @��            ����>��U?0��Cl�4          )��_�                �(��?0��        C5    T�v'&              �@  ?�  ��            "�v'&          2�  �zAd���(�          ]}��                    =���            