   �O�    ��                              �Nztv          @_��?��U���              $Nztv          @_��� �ֿ��              �Nztv          ?�����Q뿫�        ´    �Nztv          �J=r��Q뿫�        ´    LNztv          ����fc���        �4    �Nztv          ���@#����        �4    Nztv          �J=r@�뇿��        Ç    �Nztv          ?��P@�뇿��        Ç    �Nztv          ?���@���@*�B    ´  Ç    BNztv          ?���@A�@*�B    ´  Ç    �Nztv          ?���<�� @*�B    ´  Ç    �Nztv          ���<�� @*�B    ´  Ç    �Nztv          ���@�{@*=g    ´  Ç    eNztv          ���@�\u@*=g    ´  Ç  