   �l                                      �d��X       	   =�Q�                B�    wa��X       	   ��\%                ´    �i��X          >k�                 B�    �q��X          ��                  B�    �U��X          �aG�                ´    r�AF-       	   ���                      �k�AF-       	   >.{                      ��AF-          >��	                      3j�AF-          ���                      *~�AF-           �#�?(�>�              �l�AF-       	   ���    >aG�              r�AF-       	   �\'    �k�!              �X�AF-       	   >.{    >W
?              ��AF-       	   >.{    �k�!              :k�AF-          ��=r���                  �l�AF-          ��\*>�=r                  [H�AF-          >��	�u                  �&�AF-          >��	>��                