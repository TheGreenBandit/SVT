   x6�/                                      �;a2T            �3)                      �;a2T                                      �;a2T            ����                      �;a2T                                      �;a2T                                    