   �0�    z�/                              ����           �#�
��G���=q        �M    ����           �u�B�p��\'BK��@�Q��I  