   �)��    E��                              _^8x           �� ���
�.|              Y���^              @   =��G        �4    f���^              ��  =��G            