   EC�M     �+                              ��y(           �����   ?���        B�    �P���               >L��@fg        Ck    �P���               ����@fg        C�     �w           ?끿J=t?���        B�    �w           ����J=t?���        B�    �w           �:�L�J=t?���        B�    9�           �����?z�        ®    9�           �������         ®  