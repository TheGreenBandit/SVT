   ���     1�P                              5}��                                      ;Ȗ0�           ��>B�]>B�]        B�    (Ȗ0�           ?�3/>B�]>B�`        B�    *Ȗ0�           ?L��?�Q�?
>        B�    )Ȗ0�           �#��?�Q�?
>        B�    ]�v'&          @   �0(�@�  ��      ?�    ?�v'&          @!G��  A�  �      ?�    _���v           �.u?��V<#��®            b���v           ��?Ǯ�#�:®            [���v           ?�?Ǯ�#�:®            A���v           ?0��?��V<#��®            B7���                ?�Q潸Q��p            <��X       	    ���                B�    a��X       
    ���                B�    c��X           ���                B�    D��X           ���                B�    >@��            >�=q>W
>?�X��  �l        C@��            ��=r>W
>?�X��  �l        ^7���                �G�<�ز�@          