   9��?     ��                              :9��?                                A�    =9��?                                Bp    >9��?                                B�    19��?                                B�    @9��?                                C    B9��?                                C4    A9��?                                CR    C9��?                                Cp    <9��?                                C�    E9��?                                C�    G9��?                                C�    D9��?                    @��    C4  C�    M9��?                    @��    C4  C�    N9��?                    @��    C4  C�    Q9��?                    @��    C4  C�    J9��?                    @��    C4  Cp    H9��?                    @��    C4  CR    I9��?                    @��    C4  C4    U9��?                    @��    C4  C    T9��?                    @��    C4  B�    X9��?                    @��    C4  B�    ?9��?                    @��    C4  Bp    F9��?                    @��    C4  A�    O9��?                    @��    C4      