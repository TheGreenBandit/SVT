   -���                                       ���                �mp�                  0n)�           ?��?�%�S��        B���  0n)�           ?����㣾S��        B���  #0n)�           ?���.V�S��        B���  &0n)�           ?�����վS��        B���  '0n)�           ?����Ģ�S��        B���  (0n)�           ?���ȶ�S��        B���  )0n)�           ?���E/�S��        B���  $0n)�           ?���k�~�S��        B���  *0n)�           ?������S��        B���  /0n)�           ?����1#�S��        B���  00n)�           ?����dU�S��        B���  20n)�           ?L��?�%>�j��      B���  40n)�           ?L�ƽ��>�j��      B���  70n)�           ?L�ƿ.V>�j��      B���  60n)�           ?L�ƿ���>�j��      B���  0n)�           ?L�ƿ�ē>�j��      B���  90n)�           ?L���Ȯ>�j��      B���  +0n)�           ?L���E/>�j��      B���  <0n)�           ?L���k�v>�j��      B���  ;0n)�           ?L������>�j��      B���  =0n)�           ?L����x�>�j��      B���  ?0n)�           ?L�����7>�j��      B���  -0n)�           �� ?�$�S��        C�Y�  50n)�           �� ��㫾S��        C�Y�  80n)�           �� �.V	�S��        C�Y�  .0n)�           �� ���;S��        C�Y�  @0n)�           �� ��ĕ�S��        C�Y�  B0n)�           �� �ȯ�S��        C�Y�  E0n)�           �� �E/�S��        C�Y�  F0n)�           �� �k�w�S��        C�Y�  J0n)�           �� ��O�S��        C�Y�  G0n)�           �� ���8�S��        C�Y�  L0n)�           �� ��t�S��        C�Y�  M0n)�           �O\4?�%>�j��  ?�  ´   H0n)�           �O\4���>�j��  ?�  ´   I0n)�           �O\4�.V>�j��  ?�  ´   P0n)�           �O\4����>�j��  ?�  ´   O0n)�           �O\4��ē>�j��  ?�  ´   N0n)�           �O\4�Ȯ>�j��  ?�  ´   Q0n)�           �O\4�E/>�j��  ?�  ´   S0n)�           �O\4�k�v>�j��  ?�  ´   R0n)�           �O\4��O�>�j��  ?�  ´   U0n)�           �O\4���#>�j��  ?�  ´   V0n)�           �O\4���K>�j��  ?�  ´ 