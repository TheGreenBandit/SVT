   �D�     	�S                              9D:�            �.�    ?338�@      ´    :D:�            �.���?338�@      ´    ;D:�           ��п��?338�@            <D:�           >u�d���U?338�@            =D:�            ?+�>��?338�?��    B�    >D:�            ?0�վ�Q�?338�?��    B�    ?D:�            >W
P?.�?W
@�P
<    C4    @D:�            ���?.�?W
@�P
<    C4    AD:�            ���?� >�p��P
<    C4    BD:�            >u£?� >�p��P
<    C4    CD:�            �.��nr?338�@      ´    DD:�            �&fl>��?338�@  BX  ´    ED:�           >u�d��\!>aG��@            FD:�           ��� ��\!>aG��@            GD:�            ?+��aG�?338�?��    B�    HD:�            ?#�	>���?338�?���D  B�    I���^              ?��>�32        �4  