   �Z�     l`6                              %>}��               =�\*=����)          �CȖ0�           ?�  >��>�\@        B�    }@Ȗ0�           ��=p>�넽L�        B�    	Ȗ0�           ?��>�넽L�        B�    �BȖ0�           ���Q>��>�\@        B�    v/w��                ?�Q�=��4            �Bw��                >�=��4            �Aw��                ����=�G��4            �=w��            ?(��?���=R��  @�        @w��            �(��?���=�q��  ��        ���Dj       
   ��G�                B�    �
7���                    @&fe              D7���                ��36>L��              �y�e                �>�B�  ��        ?=f�M               �\(=u�B��  ´  C4    r$��Dj          �k�                 B�    _8��Dj          �k�                 B�    �4��Dj       	   ��G�                B�  