   �O�    �8o                              XK=$               �aG�>B�]        C7  