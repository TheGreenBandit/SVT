   Cw�T    =Z�                              @5ɩ4               �B�\��z�A}�        