   �     :                              ��_                    ?�              �JF��            ?\%?��>L��        ¶    G�
�                �   ?���        C7    N���v            >���=���?�fg              B���v            >L��=���?�fg              ����v            2�  =���?�fg              D���v            �L��=���?�fg              V���v            ����=���?�fg            