   9�    T�@                              }!�D�                �8Q�8Q�              ;)D:�           �u>Y?�Y�8      �4    �%D:�           >aG�>Y?�Y�8      �4    *Ȗ0�            �z�?���>��        B�    'Ȗ0�            ?̾?���>��        B�    9+�a/�            �5>�����    B�  C4    �%�a/�            ?ffR>�����    B�  C4  