   2,��                                      ����                <#�
��Q�              �%Z_�       	   �aG�                ´    �%Z_�       
   �aG�                ´    �%Z_�          �Z                ´    �%Z_�          �Z                ´    ����v           =��aG�>k�!´            ����v           >���aG�>k�!´            ����v           ?��ϾaG�>k�!´            ����v           ?����aG�>k�!´            ����v           ?�������L��´            ����v           ?�p�����B�]´            ����v           =�����B�]´            ����v           =�����#�
´          