   �As                                      	�               �fg����            