   ���                                      o~��q                   ����              u~��q              �   =L�               �l~��q              ��  =L�               �l~��q          �       =L��              �~��q          A      =L�п�            ;a~��q           ?�  �   ����        ´    �[~��q           ?�  �   ����        �4    �V~��q           ?�  �   ����        Ç  