   �$�     ��@                              <�$�                            �        h1�$�                            A�        �G͓��           ��      ��    �4       �Et_3�              A   ��          �4    <@t_3�              A�  ��          C4  