   ���     	R�                              }��                                      �Ȗ0�           ��>B�]>B�`        B�    �Ȗ0�           ?�3/>B�]>B�`        B�    �Ȗ0�           ?33(?�Q�?
>        B�    �Ȗ0�           =��s?�Q�?
>        B�    �Ȗ0�           >�̶�W
:?�         B�    �Ȗ0�           ?L̻�W
:?�         B�    �Ȗ0�           <��ʾW
:?�         B�    �^֨^           ���ƾ�(�?s3,��  �  =��	  �^֨^           ?Ǯ��(�?33 ���A�  C�
>  �^֨^           ���;�(�>�� @�Q��  B�(�  �^֨^           ?p�Ѿk�>�z�@�Q�Bx  A1G�  �^֨^           ��33���׾L�0���    B�(�  �^֨^           ?ٙ��Q�?L̴@�Q�B(  A�
P  �n�~           ��  �   ?�      ��        �n�~           ?�  �   >�
:              �n�~           �fff?� ���              �n�~           �fff����>���        �bff  �n�~            ?�  ��                    ���L                ��  ��                ���L                ��  �              