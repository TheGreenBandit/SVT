   	q��                                      �Ȗ0�            ���@   >��         B�    �Ȗ0�            ?�Y@   >��         B�    'Ȗ0�            ?��>��>�         B�    SȖ0�            ���>��>�         B�    h7���               �fg?332        B�    �@��                >��U?0��Cl�4          �@��            >���>��U?0��Cl�4          c@��            ����>��U?0��Cl�4          �
��_�                �(��?0��        C5  