   �O�                                      ��B�,       
   >�
9>��                  C	�B�,       
   >�
9=L��>B�]B�            	�B�,          >�
9=L��>B�]B�            S	�B�,          >�
9>��=��	� ��          �	�B�,          >�fa>u�Y�p� ��          �	�B�,          >�f`>u?��� ��          ��B�,          >�f`>u?��� ��          :
�B�,          ���>u>\�� ��          J
�B�,          ?���>u>\�� ��          �	�B�,       
   ?�>k����� ��          
�B�,       
   ?�>��?�f|� ��          �
�B�,       
   ����>��6]  � ��          �
�B�,       
   ?�
<>��6]  � ��        