   �O�                                      ��B�,       
   >�
9>��                  C	�B�,       
   >�
9=L��>B�]B�            	�B�,          >�
9=L��>B�]B�            S	�B�,          >�
9>��=��	� ��        