   �l     ��                              p��Dj       	                   A`  B�    ���Dj                          A`  B�    L��Dj          >�             A`  B�    6��Dj          >�            A`  B�    ���Dj          ?=p�            A`  B�    ���Dj          ?��            A`  ´    ��Dj          ��             A`  B�    ���Dj          ��            A`  B�    ���Dj          �:�A            A`  B�    ���Dj          �z�>            A`  B�    ���Dj       	   �k�             A`  B�    ���Dj       	   >aG�            A`  ´    ��8�f                ?(�?��              1�8�f                ?.z>�G�              �8�f                ??��>�\,              ��8�f                >�3<>��DB0            ��8�f                =���>��UA�            ��8�f                ��H>��T�.�          �7���            �#�
=#�
��G�A�          