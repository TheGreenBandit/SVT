   �l     1�x                              ��0�>       	                             �0�>                                    ��0�>              >���>�               ��0�>          ������Q�            