   �D�     �3                              �D:�            �.�    ?338�@      ´    OD:�            �.���?338�@      ´    �D:�           ��п��?338�@            KD:�           >u�d���U?338�@            �D:�            ?+�>��?338�?��    B�    ,	D:�            ?0�վ�Q�?338�?��    B�    �D:�            >W
P?.�?W
@�P
<    C4    D:�            ���?.�?W
@�P
<    C4    D:�            ���?� >�p��P
<    C4    2D:�            >u£?� >�p��P
<    C4    �D:�            �.��nr?338�@      ´    %D:�            �&fl>��?338�@  BX  ´    D:�           >u�d��\!>aG��@            D:�           ��� ��\!>aG��@            �D:�            ?+��aG�?338�?��    B�    @D:�            ?#�	>���?338�?���D  B�  