   �]�     >                              T}��                >B�\=�@@            OȖ0�           ��=p>���            B�    <Ȗ0�           <��'�k�=L���$  ��  B�    ����v           >� ?��Ǿ���´            ����v           =��?��Ǿ���´            X���v           ��Q�?��Ǿ���´            ����v           ���?�u����´            B7���               �B�U��Q�              ��y�e               ���    ´            �����               @�=�H    B�  B�    �%Z_�       	   ���                B�    �%Z_�       
   ���                B�    %Z_�          ���                B�    �%Z_�          ���                B�    c�V           ��Q�@G�<���A@  C4  C4    �=f�M               ��f_>�34  B�        	�V           >�@G�<���A@  C4  C4  