   �3�                                      C	����                ����L��        �4    �����                �+��L��        �4    l	�k0       	    �#�                B�    �	�k0       
    �#�                B�    \	�k0           �#�                B�    ��k0           �#�                B�  