   2,��     2
                              ����                <#�
��Q�              �%Z_�       	   �aG�                ´    x%Z_�       
   �aG�                ´    �%Z_�          �Z                ´    �%Z_�          �Z                ´    e���v           =��aG�>k�!´            ����v           >���aG�>k�!´            h���v           ?��ϾaG�>k�!´            v���v           ?����aG�>k�!´            ����v           ?�������L��´            m���v           ?�p�����B�]´            ]���v           =�����B�]´            b���v           =�����#�
´            p�v'&          =������@���C          