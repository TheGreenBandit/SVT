   ͓��     %�                              7� r           �W
D>�zᾊ=r        ¶    K� r           >��R>�zྊ=r        ¶    N� r           �aG��?����=r        ¶    H� r           >�z߿B�T��=r        ¶    j�N�"          <�                    