   �y��     .E�                              F}��            �#�
=�Q��G�              E�y��            ��                      ��Dj       	    ��                ´    "��Dj       
    ��                ´    ��Dj           �u                ´    +��Dj           �u                ´    ����v            �(�?޸T�L�´            ����v            �8Q�?�Q���'´            ����v            ��Y?����[�´            ����v            >�G�?����[�´            ����v            ?z�?޸T�L�´            ����v            ?5?�
@���'´            �Ȗ0�            ����>����բ        B�    >Ȗ0�            ?��Q>����բ        B�  