   �$�     �wj                              �F�$�                            �        GD�$�                            A�        �C͓��           ��      ��    �4     