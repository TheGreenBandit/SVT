   �O�                                      1�&O]       
   �L��        B�      ´    a�&O]          �L��        B�      ´    \�&O]          �L��        B�      ´    U�&O]       	   �L��        B�      ´    ��&O]          2�  ����>#�
        ´    ��&O]          2�  ����        B���´    ��&O]          2�  �끾�     B���´    C�&O]          �L�;�p���      B����<  7�&O]          �aG���Q�=#�    B����<  s�&O]          >u���=#�    �\
>�<  ��&O]          >�z�Ǯ��      B���ó��