   ց     _�n                              s���v            �
9?�p�>�K�´            ����v            �?��?˅">���´            ����v            ?@ 0?Ǯ?*�´            ����v            ?
9?�p�>�K�´            ]1A�           �
=m?�p�?aG�        B�    �1A�           ?�?�p�?aG�        B�    1A�           ?��>#�7?z�        B�    �1A�           ���>#�7?z�        B�    �}��                   ?
=m              ^JF��            ��z�?��?��        ´    �JF��            >W
>�?��?��        ´  