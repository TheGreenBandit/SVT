   �O�                                      <=f�M           >u>�>�fa    B�  B�    b=f�M           �k�$>�>�fa    B�  ´    =f�M           ��(��<�    ´  ´    ==f�M           <����<�    B�  ´    �=f�M           >Ǯ��<�    B�  Ç    ��8�f           ����Y��>�)              u�8�f           ����Y��?
D              �8�f           >��Y��?
D              ��8�f           >��Y��>�G�              D��Dj       	               �4      B�    h��Dj       	   �u        �4      B�    f��Dj       
   �u        �4      B�    ���Dj       
   <�        �4      B�    ��Dj          <�        �4      B�    ��Dj          ��Q�        �4      B�    #��Dj          �&fa        �4      B�    3��Dj          �&fa        �4      B�    ���Dj          �Z        �4      B�    Q��Dj          ��        �4      B�    KȖ0�           ��?xQ�?h��        B�    �Ȗ0�           =�G�?xQ�?h��        B�    Y��Dj          ����        �4      B�  