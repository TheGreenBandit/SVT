   �O�                                      &k���            �u��>.{        B�    (	k���            =�\(>�p�>.{        B�    �k���            =�G�>�Q�>.{        C�    xk���            >B�\��>.{        C�  