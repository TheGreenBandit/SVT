   @�     W                              _��3�           ��fh��3+@�              W��3�           ?�(���3+@�              R���           @
7�(Q�?�(�        C4    S���           �f`�)��?�Q�        C4    fȖ0�            ��@1G�?��        B�    UȖ0�            >���@1G�?��        B�    `����                ?L��@           C,    iP�!�               �� ?\(�        B�    e�)=�               ��  @Q�              +�z                    @�                �+�z            �\���(Q�    ´      B�    �+�z            �\����G�    ´      B�    �+�z            �\���)p�    ´      B�    �+�z            �\���
V    ´  �H  C#  