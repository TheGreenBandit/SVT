   	�%��                                      8�+            ?!G��xQ�=u              :��Dj       	    ��                ´    ;��Dj       
    ��                ´    <��Dj           @\(                B�    =��Dj           ��                ´    >��Dj       
    ��30                ´    @��Dj           @#�                B�    A��Dj           ?u                 B�    B��Dj           ?�G�                B�  