   �D�    x�c                              VH_�d               �.u>u              WH_�d               <��>u              XH_�d               >�\*=u��            YH_�d           <#�
?\&���L            ZH_�d           <#�
��G�>k�:¼      �5    [H_�d           <#�
��G�?�      �5    \H_�d           ���¿5>�3>  @*=v��    ]H_�d           ��������>�3>  @*=v��    ^H_�d           ��Q�?J=^>�(�  @*=v��    _H_�d           ���?=p���̘  @*=v    `H_�d           ���>aG���̘  A�=r    aH_�d           ����=z=�G�\<B���@    bH_�d           >B�z?�=���ª  A|Q�É    cH_�d           >B�z���=���ª  A|Q�É    dH_�d           >B�x���=u��ª  ���
É    eH_�d           >B�x�\(�>��  �&�HÉ    fH_�d           >B�x��3H>�=��k�?���É    gH_�d           >B�x?�v>�=��k�?���É  