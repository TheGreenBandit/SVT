   	�                                      ��i��                   >�Q�              b�2�           �
9���A>8Q�    ´        ��2�           �
9�f_>8Q�    ´        L�2�           ?
=n�>8Q�    B�        �2�           ?
=n�k�>8Q�    B�        G�2�           ?
=n��>8Q�    B�        ��2�           ?
=n��>8Q�    B�  ´      �2�           >�����>8Q�    B�  ´    �2�           �!G���>8Q�    B�  ´  