   �i��                                      ��                =L�о�
9              �2�           ?�M��  ���    B�        G�2�           ?�M�p����    B�        	�2�           �\,�p����    C�        ��2�           �\,��ff���    C�        f�2�           �\,�����    C�  B�    X	�2�           ?�������    C�  B�    �	�2�           ?�M�p�?L��    B�        �	�2�           ?�M���?L��    B�        �	�2�           �\,��?=p�    C�  B�    �	�2�           ?(���?=p�    C�  B�    �	�2�           �\,��ff?G�    C�        B	�2�           �\,�v?G�    C�      