   �O�     T��                              �TE$�            >k�N�W
@=�G�        ´    zTE$�            ��ֿW
@=�G�        ´    �TE$�            �B�/��=�    ´  ´     VE$�            �k��>���>.x    ®  Å    �TE$�            >k�n>�>.x�4  ¼  È�   UE$�            >W
m��=�    ´  ´     NE$�                ?��9��    �4        XUE$�                ?xQ�>lÅ  �4  C4    �UE$�                ����=�� �3  �4        7VE$�                ����?��²  �4        �UE$�            >k�N��z=�G�        ´    SUE$�            >k�N����=�G�        ´    KE$�            ��ֿ�z�=�G�        ´    �PE$�            ��ֿ���=�G�        ´    �TE$�                �#�&=��/  �  �4    �TE$�            >�z�?�(�\(@�  �4  ´    	E$�            >�z�?Y���\(@�  �4  ´    3UE$�            ���`?Y������@�  �4  B�    �TE$�            ���`?�(�\(@�
��-��B�  