   �O�     ��                              J��g-               ��\P?�XB�            .��g-               ����?(�´            /��Dj       	   �:�A                ´    H��Dj       
   �:�A                ´    G��Dj          �:�A                ´    P��Dj          �:�A                ´  