   .Å�    �u
                              �*Rf�            ��y�z྅�<��
    C7    [&�y�e           �� �p�            >��A  �*�y�e           >�=r�p�            >��A  �)�y�e           >�=r���            >��A  �+�y�e           �������            >��A