   
P�!Z                                      �� |b           ���    >��              � |b           ��ҿ���>��              d� |b           ������>��              0� |b           ����Y��>��              k� |b           ?+�    >��              �� |b           ?+����>��              E� |b           ?+��3,>��              A� |b           ?+��Z=e>��              J� |b           ?+�����>��              _� |b           ��(�����>��            