   ��m                                      �Ȗ0�          ?5 �\(�B�@�У�B�  @�    �Ȗ0�          �(ڿ^�L�8QпУ�B�  @�    �Ȗ0�          >ǮL�^�L>���B��qB�  @�    �Ȗ0�          ��Q��^�L>���B��qB�  @�    ����v           �#������L��´            ����v           ?#������L��´            ����v           >�O־���M´            ����v           ��뉾���M´            ����v           ��\.����´            ����v           >�\%����´            �%Z_�       	   �B�]                C�    �%Z_�       
   �B�]                C�    �%Z_�          ��z�                C�    �%Z_�          ��z�                C�  