   9�                                      �(�E	            ������fh>�               d(�E	           >�����fh>�               �
�E	           ��  ��fh>�             