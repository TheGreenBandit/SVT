   :��E                                      c���               �� >�AN              Ȗ0�          ����>#�
        B�    FȖ0�          =��%��>#�
        B�    "
Ȗ0�          >���?�넽��        B�    nȖ0�          ?���?����        B�    ���_�               >8Q�?���        C4  