   c"��    F�+                              �
�          ��                        ��            ?�                        q�            =���?� ?�                ��            =���@  ?���              ��            =���@&fe?�fg              e�            =���@331?�               ��            =���@?��?���              `�            =���@L��?ٙ�              r
�            =���@_��?ٙ�              ��            =���@s3-?�fh              �
�            =���@���@��            