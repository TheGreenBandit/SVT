   �#)    ���                              �����           ����    �� �        ¶    �l8�           ?   >���?
=r?333�fb      Hl8�           �#��>��?��?0����      "l8�           >���>���?
=r��f��Nf�A��  Wl8�           �   >���?
=r��f����A��