   �wb     �1                              �~�T           @�  ��  @@                �~�T           ��  ��  @@                �~�T           ��  ��  @@                �~�T           ��  ��  @@  ��      B8    �~�T           �   @@  @@          B8    �~�T           ��  AP  @@          �    �~�T           A  @�  @@          �\    �~�T           @   ��  @@                �~�T           �   ��  @@                �~�T           ��  ��  @@                �~�T           ��  ��  @�                �~�T           �   ��  @@  ��      B8    �~�T           �0  ��  @@  ��      B8    �~�T           @   @�  @@  ��      �     �~�T           ��  A  @@  ��      �   