   �$�     !=                              �t_3�           >#�
��U�7
:´          