   ���     ���                              �,}��                                      �-Ȗ0�           ��>B�]>B�]        B�    %(Ȗ0�           ?�3/>B�]>B�]        B�    s-Ȗ0�           ?33(?�Q�?
>        B�    �)Ȗ0�           =��s?�Q�?
>        B�    �+Ȗ0�           >�̶�W
:?�         B�    �-Ȗ0�           ?L̻�W
:?�         B�    #$Ȗ0�           <��ʾW
:?�         B�    6,�v'&          @   �0(�@�  ��      ?�    �-�v'&          @!G��  A�  �      ?�    -���v           �.u?��V<#��®            �%���v           ��?Ǯ�#�:®            e*���v           ?�?Ǯ�#�:®            �.���v           ?0��?��V<#��®          