   1���                                      �1���                   3   @       �4    ���Dj       	    �L��                B�    E��Dj       
    �L��                B�    7��Dj           �L��                B�    U��Dj           �L��                B�  