   �                                      �$��_                    ?�              �!JF��            ?\%?��>L��        ¶    ]'�
�                �   ?���        C7    c)���v            >���=���?�fg              �%���v            >L��=���?�fg              �(���v            2�  =���?�fg              �'���v            �L��=���?�fg              �%���v            ����=���?�fg            