   �cA�                                      �	��8                ���>��	              �	��8            ���B���>��	              ;��8            >��B���>��	              �	�J�            ��  ���E        Ç  C�    +�J�            ?� ���E        �� B�   �	��{T                @
=p>�p�    ´  C4  