   ���     L'                              ���M                                A�    6��M                                A�    8��M                                B4    ���M                                Bh    ��M                                B�    >
��M                                B�    ]��M                                B�    l��M                                B�    ~��M                                C    M��M                                C    g��M                                C    u��M                                C+    /��M                                C8    ��M                                CE    ���M                                CR    ���M                                C`    0��M                                Co    ���M                                C~    ��M                                C�    I��M                                C�    ��M                                C�    ���M                                C�    ���M                                C��   w��M                                C��   ���M                                C�� 