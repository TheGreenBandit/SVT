   ��.Q     b�V                              S1���                =�Q�=#�>���          e	���       	    ���                      ,���       
    ���                      w���           ���                      #���           ���                      ?	���       	   �Ǯ                      	���       
   �Ǯ                      h���          �Ǯ                      z���          �Ǯ                      s@��            ��p�>\?�z�        C4    �@��            ��>\?�
5        C4    o@��            =�G�>\?�
5        C4    u@��            >�p�>\?�3+        C4    �@��            ?J=p@��#��        C4    ^@��            �J=b@��#��        C4    �@��            ���U@��L��        C4    �@��            >#�&@��L��        C4  