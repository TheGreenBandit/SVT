   c"��     C�                              i|{B           A`      �Y        Cx    j|{B           A`  >8Q�A���        C�    k|{B           A`  >�=qBz�        C��   l|{B           A`  >�p�BJ�        C�    m|{B           A`  >�G�B�B�        C�    n|{B           A`  >�B�B�        C��   o|{B           A`  ?\%B�B�        C�    p|{B           A`  ?+�B�8Q        C��   q|{B           A`  ?L��C�(        C��   r|{B           A_
<?��C�(        C�    u����           A_�?���C&�>        @�  