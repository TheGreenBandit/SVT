   @�     ٪-                              �	��3�                ��  @                 M	�v�n               ��  ?B�              n	<
�            ��fe�   ?ٙ�    B�        /	<
�            ��fe�   @,��    B�        l	<
�            ��fe�  @FffB�  B�        t	<
�            ��fe�@  @FffB�  B�        �<
�            ��fe�  ?���B�  B�        �	<
�            ��fe�C37?��B�  B�        �<
�            ��fe����@*=s��  B�ff>L��  	<
�            ���	���?�z꿀  B�ff>L��  (	<
�            ��G���G�?��cB�  B�        e	<
�            ��G���=r?� B�  B�        	<
�            ���	�θR?�z꿀  B�ff>L��  �<
�            ���	�θR@*=s��  B�ff>L��  �	<
�            ���	���@*=s��  B�ff>L��  �<
�            ���	���?�z꿀  B�ff>L��  �<
�            ���	���?�z꿀  B�ff>L��  N<
�            ���	���@*=s��  B�ff>L��  ^	<
�            ���	�
��?���&  B�ff@��  �<
�            ���	��2@3��&31B�.@\,  L	<
�            ���	���N@�!�&  B�ff@��  k	<
�            ���	�.�s?�z꿀  B�ff>L��  �	<
�            ���	�.�s@*=u��  B�ff>L��  �	<
�            ��\'�#��@FffB�  B�        �	<
�            ��\'�5p�@FffB�  B�      