   �D�    %;                              ����           ?���                ���  ����           ?���?�              �>��   ���           =���?�              �>��  ���           �ffd?�      ��  @@  «34  ���           �ffd        ��  @@  «34  ����           �ffd��      ��  @@  «34  ����           =��࿀      ��  @@  «34  ����           ?��ο�      ��  @@  B	��  !���           =���    ?�  ��  @@  B	��  2���           =��࿀  ?�  ��  @@  B	��  
���           =��࿀  ?�  ��  @@  B���  �ޡ                    ?�              