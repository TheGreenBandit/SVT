   c"��                                     _B��           �O��@�����fc@�  �
33BT    4E��           �0��?�fb�W
=�'����ffB�31