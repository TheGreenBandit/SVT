   P�!Z                                      ��� P           �#�
����>�\*        ´  