   .���    �t                              Q�y�e           ���U�3���
#              w�y�e           ���U�3�>��h              ��y�e           ���U��
�>��h              U�y�e           ���U@%�>B��              a�y�e           �#���3�>���    <��
      y�y�e           ?����3�>���    <��
      �y�e           ?����&f�>���    <��
      �y�e           ?���@3.>���    <��
    