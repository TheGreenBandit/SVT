   q��     1<                              qȖ0�            ���@   >��         B�    rȖ0�            ?�Y@   >��         B�    sȖ0�            ?��>��>�         B�    tȖ0�            ���>��>�         B�    h7���               �fg?332        B�    �@��                >��U?0��Cl�4          �@��            >���>��U?0��Cl�4          c@��            ����>��U?0��Cl�4          y��_�                �(��?0��        C5    m�v'&              �@  ?�  ��            }�v'&          2�  �zAd���(�        