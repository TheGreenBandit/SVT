   �D�    2�                              �H_�d               �.u>u              �H_�d               <��>u              �H_�d               >�\*=u��            �H_�d           <#�
?\&���L            �H_�d           <#�
��G�>k�:¼      �5    �H_�d           <#�
��G�?�      �5    �H_�d           ���¿5>�3>  @*=v��    �H_�d           ��������>�3>  @*=v��    �H_�d           ��Q�?J=^>�(�  @*=v��    �H_�d           ���?=p���̘  @*=v    �H_�d           ���>aG���̘  A�=r    �H_�d           ����=z=�G�\<B���@    �H_�d           >B�z?�=���ª  A|Q�É    �H_�d           >B�z���=���ª  A|Q�É    �H_�d           >B�x���=u��ª  ���
É    �H_�d           >B�x�\(�>��  �&�HÉ    �H_�d           >B�x��3H>�=��k�?���É    �H_�d           >B�x?�v>�=��k�?���É    ^t_3�          >B�]�  �^�P®          