   v*�    P�5                              "v*�                           �         �v*�                           A         �v*�                           A�        ?v*�                           ��        Uv*�                           �H        �v*�                           BH      