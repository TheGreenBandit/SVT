   c"��     )�O                              ��           ��                        �           ?�                        ��            ���T?�38>��Q              ��            �\,@  ?\(�              ��            =��@&fe?�fg              ��            �#�J@331?�               ��            <#��@?��?�z�              ��            =���@L��?�G�              ��            =���@_��?�
>              ��            =���@s3-?�fh              �            =���@���@��              �                @�  @$z�            