   	����     �D                              ��J�            ?   ��    ����          ��J�            �   ����    �噘=���      �J�            �.y���    ��            ��J�            >#�
����    �陖          *��8            �  ���?�fb    C4        ���8            �  ���?�fb    C4        ���8            ?����?�fc    C4        ��{T            >���?332?˅��\(B�3;�1��  ��{T            ���?.z?˅��\(B�3;�1��