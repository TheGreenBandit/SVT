   �O�     9Zn                              �GY^&                �ٙ�����              �GY^&                ?�  ����              �%Z_�       	    @~                ´    �%Z_�       
    @~                ´    �%Z_�           @~                ´    �%Z_�           @~                ´    ����^              @�              C4    ����^              ��G�@&fdA      C4  