   ��     4�                              "͓��                            C4        <o���            ?�fg    ���?�  ��      	o���            ����    ���?�  B�        �V            ��Q�?334                  t�V            �
=���=���              ^�V            >W
>���=���              R�V            >W
>��¾���              ��V            ���G��¾���              #�y�e                �33<�´            E�y�e            �����>�z�´            z�y�e            ����̾aG�´            S�y�e            >B�\��̾aG�´          