   
�]�     �Z�                              5�]�           �334                      6}��               =���=�����            7}��           �:�L=�Q�=�����            8Ȗ0�           ��Q�@ ��>L��        B�    9Ȗ0�           �\(�@ ��>L��        B�    :Ȗ0�           >u@ ��>L��        B�    ;Ȗ0�           ��fg>W
&58          B�    <Ȗ0�           ?��>W
&58          B�    BJF��               ����>�\)        ³ǫ  CJF��           �J=t����>�\)        ³ǫ