   {~V�                                      �{~V�           @�                        �{~V�            @�  �@��@p�´            {{~V�            @�  �@��@���´            w{~V�            @@  �@��AQ�    ²  ´    ]{~V�                �@��@p�´            �{~V�                �@��@�Q�´            y{~V�            @���@��A<��´            A{~V�            @���@��Ap)´            �{~V�            �����@��A�z�    �4  B�    i{~V�            @����@��A�z�    �4  C�    �{~V�            @���@��A��B�      C4  