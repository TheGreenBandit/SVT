   ��    B��                              Qp��                    ?�                4Qp��            >���    ?�                ZQp��            �      ?�                �Qp��            �ffh    ?332              �Qp��            ?ffg    ?332              .Qp��            ?ffg    >���              FQp��            �ffh    >���              Qp��            ����    ?�34              $Qp��            >���    ?�34              �Qp��            ��      ?ٙ�              TQp��            ��  @��@l���   �   ®    WQp��            ��  @��@,��´  ��  ®    �Qp��            ��  @��@l��´  ��  ®  