   /T{    3�W                              D	�               >�z�?Tz�            