   ͓��     6�                              �� r           �W
D>�zᾊ=r        ¶    �� r           >��R>�zྊ=r        ¶    �� r           �aG��?����=r        ¶    �� r           >�z߿B�T��=r        ¶    ��v�n          ��G�                      #�v�n          ?�\'                      ����^              AC�"���        �4    ����^              A�?��@�      �4  