   	�O�    3Q                              
�8�Q                                �     h	�8�Q                                º    �	�8�Q                                �4    "	�8�Q                                Æ    �	�8�Q                        B(  ��  �4    �8�Q                        C  �I  �4    ^	�8�Q                        C;  �7  �4    _	���^              @@              C4    g	���^              �@                  