   c"��     �z                              #|{B           A`      �Y        Cx    $|{B           A`  >8Q�A���        C�    %|{B           A`  >�=qBz�        C��   &|{B           A`  >�p�BJ�        C�    '����           A`      B�          ��  