    ���                                      ��γ�           ��fh    ��          ´    �γ�           ��fh    ��      ��  ´fh  <�γ�           ?�fe    ��  �4  ��  ´fh  O%�γ�           ?�fe    ��  �4  �q��¶��  6$�γ�       	    ?�fe    ��  �4  �q��¶ff  �&�γ�       	    ?�fe    ��  �4  �#��¶ff  G�γ�       	    ��fl    ��  ô  ���¶ff  	�γ�       	    ��fl    ��  ô  ����¶ff  ��γ�                    >L���%           w$�γ�            =���    >L���%           ��γ�            ����    >L���%           ��γ�            ����    =����%           �!�γ�            ��      =����%           �/�γ�            =���    =����%           �#�γ�            =���    2�  �%           �9�γ�            ��      2�  �%           �"�γ�            ����    2�  �%         