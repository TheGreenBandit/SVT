   E�j�                                      �E�j�                                C4  