   �$�     �(                              �E�$�                            �        n/�$�                            A�        �>͓��           ��      ��    �4       �Ht_3�              A   ��          �4    q0t_3�              A�  ��          C4  