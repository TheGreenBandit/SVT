   �     �B                              &D:�            �O\,�\(�?��        ²    3D:�            �O\,��(�?��        ²    AD:�            �O\,�z�?��        ²    aD:�            ���X���?��              OD:�            �������?��              DD:�            >��s���?��              �D:�            ?L̺��?��        B�    D:�            ?L̺�T?��        B�    )D:�            ?L̺�k�?��        B�    bD:�            >��,�\(?��        C4    YD:�            �0  �\(?��        C4    5D:�            �  �\(?��        C4  