   �$�     ��                               @o�$�                           �        �i�$�                           A�        �l͓��           ��      ��    �4       7it_3�              A   ��          �4    ct_3�              A�  ��          C4    Ctt_3�              A�  ��          C4    wst_3�              A�  ��          C4    $`t_3�              A�  ��          C4    e_t_3�              A   ��          �4    �kt_3�              A   ��          �4    	Xt_3�              A   ��          �4  