   ͓��                                      R� ��       	    ?�G�            ´        <� ��       
    ?�G�            ´        e� ��           ?�G�            ´        ]� ��           ?�G�            ´        y� ��           <#�*�(����p�              a� ��           <#�*��  ��p�              }� ��           <#�*?z��y��            � ��           <#�*��)��=t¬            6� ��           <#�*��(��33H¬      C4    K� ��           ��3*�\(`�z�´      C�    >� ��           ��3*�,̠��,´      C�    �� ��           ��3*?aH2�� ´      C�     � ��           ?�Q��,̠�z�´      B�    Y� ��           ?�Q��Y��z�´      B�    z� ��           ?�Q�?G�����N´      B�  