   KlV�     Z�                              U7���            2�      ?�fh              V7���            ����L��>L���f�          W7���            2�  ?   ?�fh              X7���           ����?   ?�fh              Y7���           >���?   ?�fh              Z7���            ?���L��>L���f�        