   �$�                                      0&��           �ff]��^?Y��B�            �&��           ?k���^?Y��B�            �
&��       	   �u�:�#�*<��WB�      B�    &��       
   �u�:�#�*<��WB�      B�    �
&��          �#׾��  �  B�
L    B�    �&��          �#׾��  �  B�
L    B�  