   	�a&                                      5��X       	   �\'        ��  �� B���  R��X       
   �\'        ��  �� B���   ��X          �W
;        ��  �� B���  D��X          �L��        ��  �� B���  'WTr�       	   �\"                ³��  QWTr�       
   �\"                ³��  SWTr�          �W
5                ³��  :WTr�          �W
5                ³��  jc"��                   >���            