   ��.Q     ��                              �
1���                =�Q�=L��>���          �
���       	    <#�                      �Oʥ            �J=i@
=q���b    B�  B�    �Oʥ            ?O\2@
=q���b    B�  B�    �Oʥ            >\J@
=q�#ն    B�  B�    �Oʥ            �\@
=q�#ն    B�  B�    ����^              @s30��        C4    :���^              ����@�@���    C4    3���       
    <#�                      j���           <#�                      !���           <#�                      M���       	   ���Q                      ����       
   ���Q                      g���          ���Q                      S���          ���Q                      ����          ���Q                    