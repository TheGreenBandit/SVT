   KlV�                                      HKlV�                        �0  =�� ��    IKlV�                        ��  =�� ��    JKlV�                        �  =�� ��    MKlV�                        �<  =�� ��    NKlV�                        �p  =�� ��    OKlV�                          =�� ��    PKlV�                        ¸  =�� ��    TKlV�                        ��  =�� ��    UKlV�                        ��  =�� ��    XKlV�                        �  =�� ��    YKlV�                        �  =�� ��    hKlV�                        �)  =�� ��    iKlV�                        �4  =�� ��    lKlV�                        �?  =�� ��    mKlV�                        �J  =�� ��    tKlV�                        �W  =�� ��    uKlV�                        �c  =�� ��    xKlV�                        �o  =�� ��    yKlV�                        �{  =�� ��    |KlV�                        Ã  =�� ��    }KlV�                        Ç� =�� ��    �KlV�                        Ë� =�� ��    �KlV�                        Ð  =�� ��    �KlV�                        Ó  =�� ��    �KlV�                        Ö� =�� ��    �KlV�                        Ú� =�� ��    �KlV�                        Þ  =�� ��    �KlV�                        â� =�� ��    �KlV�                        è  =�� ��    �KlV�                        í� =�� ��  