   ͓��                                      )`��G       	    ��d                C�    !`��G       
    ��d                C�    %`��G           ��d                C�    p`��G           ��d                C�    �`��G       	    �p                C�    B`��G       	    �aG�                C�    `��G       	    �#׾                C�    E`��G       	   >#��                C�    ``��G       	   >�c                C�    f`��G       
    �p                C�    `��G           �p                C�    g`��G           �p                C�    ~`��G       
    �aG�                C�    �`��G           �aG�                C�    �`��G           �aG�                C�    �`��G       
    �aG�                C�    �`��G           �aG�                C�    x`��G           �aG�                C�    �`��G       
    �#׾                C�    �`��G           �#׾                C�    �`��G           �#׾                C�    �`��G       
   >#��                C�    �`��G          >#��                C�    �`��G          >#��                C�    w`��G       
   >�c                C�    #`��G          >�c                C�    `��G          >�c                C�  