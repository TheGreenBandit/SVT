   ���     �r�                              �}��                                      �Ȗ0�           ��>B�]>B�]        B�    �Ȗ0�           ?�3/>B�]>B�`        B�    �Ȗ0�           ?L��?�Q�?
>        B�    �Ȗ0�           �#��?�Q�?
>        B�    ��v'&          @   �0(�@�  ��      ?�    ��v'&          @!G��  A�  �      ?�    ����v           �.u?��V<#��®            ����v           ��?Ǯ�#�:®            ����v           ?�?Ǯ�#�:®            6���v           ?0��?��V<#��®            �7���                ?�Q潸Q��p            ���X       	    ���                B�    ���X       
    ���                B�    b��X           ���                B�    ���X           ���                B�    �@��            >�=q>W
>?�X��  �l        �@��            ��=r>W
>?�X��  �l        �7���                �G�<�ز�@            ��y�e                ��_    ´            �w��                    B�  �4          