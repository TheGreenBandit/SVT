   �%��                                      @$                ��G���Y              ���Dj       
                       ´    {��Dj       
   �L��                ´    ���Dj                              ´    ~��Dj                              ´    ���Dj                              ´    -��Dj          �L��                ´    ���Dj          �L��                ´    ���Dj       	                       ´    F��Dj       	   �L��                ´    N�l�                ?�\!=�H<��
    C4  