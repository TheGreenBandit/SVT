   
�]�     EU                              �M}��                >B�\=�@@            Ku�v'&              ����@��KC            �mȖ0�           ��=p>���            B�    �uȖ0�           <��'�k�=L���$  ��  B�    �>���v           >� ?��Ǿ���´            �n���v           =��?��Ǿ���´            ����v           ��Q�?��Ǿ���´            X=���v           ���?�u����´            �D7���               �B�U��Q�              P�y�e               ���    ´          