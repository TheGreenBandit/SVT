   �#)                                     +��	�               ����>L��=#�
<#�
C/  