   ��                                      ^�V            >���?       ����          c�V            �� ?\(�#�
@�R�����4�Z  _�a/�            ��Q�>�>�\(B�  ´��B�ff  e�a/�            ��Q�?(��>�\(B�  ´��B�ff  g�a/�            ��p�?^�O>�\(B�  ´��B�ff  i�a/�            ��p�?^�O>�\(B�  ´��B�ff  j�a/�            >��e?^�O>uB�  ´��¯��  l�a/�            >��e?#�>��B�  ´��¯��  �a/�            >�̭>���>uB�  ´��¯��  (�k0       
                        µ��  !�k0       	                        µ��   ��Dj                               ´    *��Dj                               ´  