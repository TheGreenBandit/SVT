   �i�    h�                              ��i�           @�                        2�i�           A                         � �i�           A       @@                ��i�                   @@                ��i�           @�      @@              