   ͓��     ��                              8`��G       	    ��d                C�    9`��G       
    ��d                C�    :`��G           ��d                C�    ;`��G           ��d                C�    <`��G       	    �p                C�    =`��G       	    �aG�                C�    >`��G       	    �#׾                C�    ?`��G       	   >#��                C�    @`��G       	   >�c                C�    A`��G       
    �p                C�    B`��G           �p                C�    C`��G           �p                C�    D`��G       
    �aG�                C�    E`��G           �aG�                C�    F`��G           �aG�                C�    G`��G       
    �aG�                C�    H`��G           �aG�                C�    I`��G           �aG�                C�    J`��G       
    �#׾                C�    K`��G           �#׾                C�    L`��G           �#׾                C�    M`��G       
   >#��                C�    N`��G          >#��                C�    O`��G          >#��                C�    P`��G       
   >�c                C�    Q`��G          >�c                C�    R`��G          >�c                C�    \o���                �� =���              ]o���            ?Tzο� ?���    ´        ^o���            �+�E�� ?���C/  B�      