   9��?    �")                              T�l��           >�=q@P��>��            