   9�                                      �D�                ����                  �D�                                      �D�                ����                  fD:�            �L��>���?L���8      C4    �D:�            >L��>���?L���8      C4    jD:�           ����>L�ξk�    B�  C�   �D:�           ?�|>L�ξu    B�  C� 