   �wb                                      8�wb                            ��        ?�wb                            A�        B�wb                            �         F�wb                            B         J�wb                            �p        O�wb                            Bp      