   
/T{    �t\                              �
-�b/           ��fa>� ���              �JF��           >��ɿ�>aG�        ²    �
JF��           �!G���>aG�        ²    kJF��           �!G���Q?�        ²    �JF��           >�p���Q?�        ²    yJF��           >�fd��3+�#��¨  ?�  ²    �JF��           >�fd��3+�#��¨  ?�  ²    XJF��           ?(����3+�#��¨  ?�  ²    ^JF��           ��Q쿳3,�#��Ç� ?�  ²    �JF��           ��Z��3,�#��Ç� ?�  ²  