   ���     (�E                              ����               �J�G                  sD:�            ?xQ�    >�=���      B�    �D:�            ?xQ�(�>�=���      B�    �D:�            ?xQ쿚�A>�=���      B�    �D:�            ?xQ����>�=���      B�    D:�            ?xQ���>�=���      B�    pD:�            ?xQ��B�R>�=���      B�    �D:�            ?xQ��h��>�=���      B�    �D:�            �p���h��>�=���      ´    D:�            �p���A�{>�=���      ´    oD:�            �p����>�=���      ´    �D:�            �p���>�=���      ´    �D:�            �p�迟��>�=���      ´    �D:�            �p��#�>�=���      ´    #D:�            �p��u��>�=���      ´    �%Z_�       	    �L��                ´    �%Z_�       
    �L��                ´    �%Z_�           �L��                ´    �%Z_�           �L��                ´    �%Z_�           �\(����G�        ´    �%Z_�           �\(��(�G�        ´    n%Z_�           ?\(���\#�M        B�    �%Z_�           ?\(���\;�M        B�    D:�            �p�����>�=���      ´    D:�            �p����Q�>�=���      ´    D:�            ?xQ����>�=���      B�    wD:�            ?xQ����?>�=���      B�  