   ��     D%�                              ;Qp��                    ?�                �Qp��            >���    ?�                QQp��            �      ?�                Qp��            �ffh    ?332              MQp��            ?ffg    ?332              Qp��            ?ffg    >���              �Qp��            �ffh    >���              �Qp��            ����    ?�34              �Qp��            >���    ?�34              PQp��            ��      ?ٙ�              Qp��            ��  @��@l���   �   ®    �Qp��            ��  @��@,��´  ��  ®    
Qp��            ��  @��@l��´  ��  ®  