   
�%��                                      
�2�               ��                  <�2�               ?z�                  `��Dj       	                       ´    ���Dj       	   �u                ´    ���Dj       
                       ´    d��Dj                              ´    ���Dj                              ´    ���Dj       
   �u                ´    ��Dj          �u                ´    ���Dj          �u                ´  