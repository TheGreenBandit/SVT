   !��}     P�0                              /!��}               ���<#�
        �4    ��B�,       
   �                   B�    �B�,          �                   B�    j�B�,          �                   B�    Z�B�,       	   �                   B�    ��B�,          �� �334�          B�    ��B�,       	   �� ��  3�          B�    }�B�,       	   @?����  3�          B�    ��B�,          @?����  3�          B�    J�B�,          @?����  3�          B�    �B�,          �� ��ff�          B�    ��B�,          @   ��ff�          B�    ��B�,          @   �330�          B�     �)=�                   @,��        �4  