   q��                                      �
 �3�            A`  �   BV��    ´        �
 �3�            A`  A  BV��    ´         �3�            @�  A  BV��    ´         �3�            @�  �   BV��    ´      