   2,��     ś�                              2f����                =��q    @             �^���            <s=�Q�q��               f��;#       	    ��                 ´    td��;#       
    ��                 ´    -d��;#           ��                 ´    Xe��;#           ��                 ´    �f���v            ?+�?�|<��
´            �e���v            ?
=s?��H<#�
´             e���v            �
=n?��H<#�
´            �f���v            �.v?���<�´            _b���v            �33.?�
>���´            cd���v            �
:?�
>���Q´            �d���v            ?��?�
>���Q´            &���v            ?33,?�
>�� ´            �\����            <#�
@=p�#�    B�  B�    �`����           �h��?�3-�33-    ��        De����           ?fft?�3-�33-    ��  C4  