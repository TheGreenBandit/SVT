   ��\�                                      �.�                =�Q�=���              ���Dj       	   �u                ´    ���Dj       
   �u                ´    ���Dj                              ´    b��Dj          ?��                ´    ���Dj          ?��                ´    ���Dj          �
9                ´    ���Dj          �
9                ´    �O{Q�               @G�=u�BB,      C4    �O{Q�           ��� @G�=u�BB,      C4    �O{Q�           >�z�@G�=u�BB,      C4    2�5�V            �ff]�}p��L��        B�    ��5�V            �ff]�}p��z�        B�    \�5�V            ?ff]�}p��z�        B�    ��5�V            ?ff]�}p��^�I        B�  