   �]�     ���                              ��]�                                �p    ��]�                                ��    S�]�                                �4     �]�                                �p    %�]�                                    1�]�                                ´    >�]�                                ��    {�]�                                ��    C�]�                                �    e�]�                                �    R�]�                                �     ��]�                                �/    �]�                                �>    h�]�                                �M    /�]�                                �\    ��]�                                �k    Q�]�                                �z    ��]�                                Ä�   E�]�                                Ì    ��]�                                Ó�   d�]�                                Û    ��]�                                â�   ��]�                                ê    �]�                                ñ�   ��]�                                ù    u���%              �ٙ�@334C          