   �y��                                     �ꕭ0            �d  BT  C�  �H  B�  B�    �ꕭ0            �x  BI=�C�� �X  B�  B�    �ꕭ0            ��  BpNC���X  B�  B�  