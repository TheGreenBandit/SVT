   �$�     �΃                              �G�$�                            �        �/�$�                            A�        �͓��           ?��    �#�&    �4       ;A͓��           �Ǯ    ���    �4        �Cl�m                ?�                  