   �O�    U�H                              �	BjT|                   >�fb        C4�