   C*�f                                      �D�                    =���              {�7                                      {�7                                      Z7���                                      Z7���                                      a<CN                ��37>���B:��          m�܇                  ��                t�܇                  ��              