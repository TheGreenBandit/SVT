   c"��                                     -3�g�@                   A`              