   1���                                      �
����                ���Z�             �
�E	            �J=i?����´            �E	            ?J=?�=z��´            �E	            >B��?�=z���´            ]�E	            �L�u?�=z���´            \�k0       	   ���                B�    ^�k0       
   ���                B�    �
�k0          ���                B�    �
�k0          ��z�                C�    =�k0          ��z�                C�    =f�M            �n|��t��բ        ´    =f�M            �n|���P��բ        ´    H=f�M            �n|��X��բ        ´    =f�M            ?h�Ŀ�t��բ        B�    =f�M            ?k� ��G���բ        B�    %=f�M            ?k� �(�ȼ�բ        B�  