   c"��                                       ���                    @�  B�            � ���                    A�  B�            � ���            A�      @�  B�            � ���            ��      @�  B�            ? ���            ��      A�  B�            � ���            B      A�  B�          