   !��}                                      �!��}               ���<#�
        �4    �#�B�,       
   �                   B�    �&�B�,          �                   B�    |$�B�,          �                   B�    g$�B�,       	   �                   B�    ��B�,          �� �334�          B�    ��B�,       	   �� ��  3�          B�    1'�B�,       	   @?����  3�          B�    )%�B�,          @?����  3�          B�    �"�B�,          @?����  3�          B�    @&�B�,          �� ��ff�          B�    �'�B�,          @   ��ff�          B�    ~!�B�,          @   �330�          B�  