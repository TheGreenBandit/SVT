   	���     Y�c                              6
}��                                      �	Ȗ0�           ��>B�]>B�]        B�    
Ȗ0�           ?�3/>B�]>B�]        B�    �
Ȗ0�           ?33(?�Q�?
>        B�    o
Ȗ0�           =��s?�Q�?
>        B�    d
�~h�            ?��                      �	~��q            �L��                      �	~��q                                      �	~��q                    ??��            