   �)��    S��                              �Fk�9           >���L�Ϳ&fa        C6  