   �O�                                      �`G�
                   �.z        �4    ��;#       	    ��<#�
���
        ´    ���;#       
    ��<#�
���
        ´    ���;#           ��<#�
���
        ´    "��;#           ��<#�
���         ´    M`G�
               ��
$��        ô    ��
�                ��p�?��
°            �
�            �W
?��p�?E�°            f�
�            >aG���p�?E�°            �Oʥ                ��h?)    �4        �Oʥ                ?B�`>�)     �4      