   �%��                                      @$                ��G���Y              �@���                �g��
9              ���Dj       
                       ´    {��Dj       
   �L��                ´    ���Dj                              ´    ~��Dj                              ´    ���Dj                              ´    -��Dj          �L��                ´    ���Dj          �L��                ´    ���Dj       	                       ´    F��Dj       	   �L��                ´  