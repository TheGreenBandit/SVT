   @�     �:[                              �!               ��p�?z�        B�  %B�<           >�(�    @           C��   ��!               ��p�@6fd        B�  a�!               ��p�@tz�        B�