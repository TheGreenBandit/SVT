   vqd�    ��                              ,}��                =�G�<#�
              }%Z_�       	   ���                B�    �%Z_�       
   ���                B�    �%Z_�          �k�                 B�    X%Z_�          �k�                 B�    +j�&�           �xQ�    �
=m        Ç    �j�&�           ?z�H    �
=m        Ç    :����                @�ֽL��    Ì  B�    ;����            >k�!@�ֽL��    Ì  B�    Y����            �� @�ֽL��    Ì  B�    ����v            �5?��L�L��´            ����v            ��?��L����´            ����v            ?�z?��L����´            <���v            ?33&?��L�L��´            �V���                �G�=�G�              s=f�M                ��35>��
3!B�      