   �(8                                      {�2�            ����?��Ծ�               ��2�            >�z�?��Ծ�=q              ��2�            ��=q>�� ���              ��2�            ��=q�Tzξ��              ��2�            ��=q��fW��z�              ��2�            >�=r��fW��\*              ��2�            >�=r��̴���              ��2�            >�=r>�����              �%Z_�       	   ����                ´    �%Z_�       
   ����                ´    �%Z_�          ����                ´    �%Z_�          ����                ´  