   
c"��    S��                              v|{B           A`      �Y        Cx    .|{B           A`  >8Q�A���        C�    ^|{B           A`  >�=qBz�        C��   x|{B           A`  >�p�BJ�        C�    t|{B           A`  >�G�B�B�        C�    n|{B           A`  >�B�B�        C��   Y|{B           A`  ?\%B�B�        C�    <|{B           A`  ?+�B�8Q        C��   X|{B           A`  ?L��C�(        C��   q|{B           A_
<?��C�(        C�  