   �O�     $��                              �8��               �����Q        ´    ���Dj       	   ����                ´    ���Dj       
   ����                ´    ���Dj          ����                ´    ���Dj          ����                ´    W��9�               ����?J=���            �{��
                ����#��            RL��<              @�              C4    QL��<              ��                    �y���            �5      A�  �4            Oy���            C�      A�  �4          