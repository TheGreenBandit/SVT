   @�     2W                              
@�           @                        ��3�           �332��  @              ��3�           @1G���  @              �.���           ?�  �Ф ?���              ��o�           ��
5�A�?aG�        B�    c�o�           >#��A�?aG�        B�    b�o�           ?�G��A�?aG�        B�    ��o�           @W
9�A�?aG�        B�    JF��           ������=?^�T        ´    �JF��           @p�����=?^�T        ´    d����            �Ǯ����?�        C4    �����            @ffh����?�        C4    �.���            ��z˿���?aG�        B�    %.���            @�Q쿿��?aG�        B�  