   (c"��     T��                              �|{B           A`      �Y        Cx    �
|{B           A`  >8Q�A���        C�    �	|{B           A`  >�=qBz�        C��   �|{B           A`  >�p�BJ�        C�    ]|{B           A`  >�G�B�B�        C�    L|{B           A`  >�B�B�        C��   �
|{B           A`  ?\%B�B�        C�    �|{B           A`  ?+�B�8Q        C��   
|{B           A`  ?L��C�(        C��   �
|{B           A_
<?��C�(        C�    S|{B           A]G�?��C)�(        CԀ   �|{B           AZ=h?��C:�(        C܀   a
|{B           AW�?��CK��        C�    |{B           AW�?k�C\��        C�    u|{B           AW�?J=jCm��        C�    ^|{B           AW
0?33.C~��        D     �|{B           AW
0?��C��        D    �|{B           AY�|?�ZC�j8        D	@   |{B           A]G�?�ZC��8        D�   <|{B           A_\(?!G�C�k�        D@   �|{B           Ac38?(��C��        D�   4|{B           Ae�?(��C�k�        D    �|{B           Ah��?(��C���        D @   p|{B           Ah)?E�C�~�        D$�   |{B           Ah)?h��C��p        D)    �	|{B           Ah)?�\#Cԅ         D-@   �	|{B           Ah)?ǮC�         D1@   v	|{B           Ah)?���C��        D5@   
|{B           Ab=t?��;C��        D9�   �	|{B           A_\(?��;C���        D=�   i|{B           A[�?��;C��        DB@   
|{B           AW��?��;D��        DF�   m|{B           AT��?�=eD�        DK�   �|{B           AT��?˅DH�        DP@   �|{B           AT��?�3+D��        DT@   �|{B           AT̼?��AD��        DX�   9|{B           AT̼?h��D�        D]    �|{B           AW��?h��DH�        Da@   s|{B           A[
6?h��D!��    ��  Df    �|{B           A`(�?z�>D%��    ��  Dj@ 