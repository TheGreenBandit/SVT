   	�Z�     '�k                              �}��               =�G�>8Q�@]p~          �Ȗ0�           ?�  >��>�\@        B�    ZȖ0�           ��=p>�넽L�        B�    Ȗ0�           ?��>�넽L�        B�    Ȗ0�           ���Q>��>�\@        B�    I��Dj       
   ��=q                ´    ���Dj          ��=q                ´    ��Dj          ��=q                ´    a��Dj       	   ��=q                ´  