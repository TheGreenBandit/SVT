   �#)                                      ~�k0       	    ��\(                ´    ��k0       
    ��\(                ´    ��k0           ��\(                ´    ��k0           ��\(                ´    p^a�                                      p^a�                                      p^a�                                      �1A�                                      �1A�                                      �1A�                                      �Rf�                ����=���        �4  