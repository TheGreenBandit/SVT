   �O�    9i                              :Nztv           @_��?��U���              �Nztv           @_��� �ֿ��               Nztv           ?�����Q뿫�        ´    iNztv           �J=r��Q뿫�        ´    Nztv           ����fc���        �4    WNztv           ���@#����        �4    �Nztv           �J=r@�뇿��        Ç    [Nztv           ?��P@�뇿��        Ç    ZNztv           ?���@���@*�B    ´  Ç    �Nztv           ?���@A�@*�B    ´  Ç    �Nztv           ?���<�� @*�B    ´  Ç    �Nztv           ���<�� @*�B    ´  Ç    �Nztv           ���@�{@*=g    ´  Ç    �Nztv           ���@�\u@*=g    ´  Ç  