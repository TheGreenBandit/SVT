   � L�                                      p �3�            Bx  �  ��                � �3�            Bx  ��  ��                � �3�            Bx  ��  ��                � �3�            Bx  @�  ��                � �3�            A0  B�  ��          B�    � �3�            �x  A�  �0  ��      C1    � �3�            �|  A   �0  ��      C3    � �3�            �|  �  �0  ��      C3    � �3�            �|  ��  �0  ��      C3    �$vM            B  A�  ��  ®            �$vM            A�    ��  ¦      ��    �$vM            ��  A�  �p  ´      B�    #$vM            �L  ����p  ´      C7fd  K$vM              �Z��B0  �@  @L��C>fd  �$vM              �Z����      �5��C>fd