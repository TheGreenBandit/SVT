   c"��     %�                              |{B           A`      �Y        Cx    |{B           A`  >8Q�A���        C�    
|{B           A`  >�=qBz�        C��   |{B           A`  >�p�BJ�        C�    |{B           A`  >�G�B�B�        C�    |{B           A`  >�B�B�        C��   |{B           A`  ?\%B�B�        C�    |{B           A`  ?+�B�8Q        C��   |{B           A`  ?L��C�(        C��   |{B           A_
<?��C�(        C�    |{B           A]G�?��C)�(        CԀ   |{B           AZ=h?��C:�(        C܀   |{B           AW�?��CK��        C�    |{B           AW�?k�C\��        C�    |{B           AW�?J=jCm��        C�    |{B           AW
0?33.C~��        D     |{B           AW
0?��C��        D    |{B           AY�|?�ZC�j8        D	@   |{B           A]G�?�ZC��8        D�   |{B           A_\(?!G�C�k�        D@   ����           A[�?!G�C��h        C;  