   c"��    .��                              $
'\                ��  B  B�            G
'\            ��  ��  B  B�            `	'\            A�  ��  B  B�            �
���%              @�  ?���C          