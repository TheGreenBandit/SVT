   �Kw�    R9�                              ��E\           ��z�n�@�        ´��