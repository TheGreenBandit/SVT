   	q��     
��                              ;Ȗ0�            ���@   >��         B�    =Ȗ0�            ?�Y@   >��         B�    Ȗ0�            ?��>��>�         B�    BȖ0�            ���>��>�         B�    !7���               �fg?332        B�    5@��                >��U?0��Cl�4          9@��            >���>��U?0��Cl�4          <@��            ����>��U?0��Cl�4          >��_�                �(��?0��        C5  