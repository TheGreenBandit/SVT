   q��     Q�                              �Ȗ0�            ���@   >��         B�    �Ȗ0�            ?�Y@   >��         B�    �Ȗ0�            ?��>��>�         B�    �Ȗ0�            ���>��>�         B�    �7���               �fg?332        B�    �@��                >��U?0��Cl�4          �@��            >���>��U?0��Cl�4          �@��            ����>��U?0��Cl�4          ���_�                �(��?0��        C5    ��v'&              �@  ?�  ��            ��v'&          2�  �zAd���(�          �}��                    =���            