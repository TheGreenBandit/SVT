   c"��                                     +�)YO            @   �A��    ´  Â    -�)YO            ��  @��A��    ´  ô    3�)YO            AJf^@��A��    ´  �	    4�)YO            ��35A#\(A+�        ��   .�)YO            ���^A(�A+�        �� 