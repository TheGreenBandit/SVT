   ���     p�~                              �	}��                    =��	               Ȗ0�           �
D?��>aG�        B�    �Ȗ0�           ?\"?��>aG�        B�    V@��           ��z@Q�W
        C4    �@��           >��	@Q�L̡        C4    �@��           �#�@Q�W
        C4    4=f�M                ��Q�>�����B�      