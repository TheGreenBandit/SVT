   	���     &!                              y}��                                      zȖ0�           ��>B�]>B�]        B�    {Ȗ0�           ?�3/>B�]>B�]        B�    |Ȗ0�           ?33(?�Q�?
>        B�    }Ȗ0�           =��s?�Q�?
>        B�    ~�~h�            ?��                      ~��q            �L��                      �~��q                                     �~��q                   @Nw            