   vqd�                                      �}��                =�G�<#�
              �%Z_�       	   ���                B�    �%Z_�       
   ���                B�    �%Z_�          �k�                 B�    �%Z_�          �k�                 B�    �j�&�           �xQ�    �
=m        Ç    �j�&�           ?z�H    �
=m        Ç    D����                @�ֽL��    Ì  B�    :����            >k�!@�ֽL��    Ì  B�    �����            �� @�ֽL��    Ì  B�    i���v            �5?��L�L��´            Q���v            ��?��L����´            ����v            ?�z?��L����´            ����v            ?33&?��L�L��´            �V���                �G�=�G�              �=f�M                ��35>���3!B�      