   �0�    |d                              �7���                <��
>�=qA��          �7���                ���A>�=q���334      �7���                                      ���I                   ��=p            