   �D�   u_                              �\��               ���	��G�        C3)