   �O�     %��                              ���Dj       	               �4  �X  B�    �
��Dj       
               �4  �X  B�    |��Dj                      �4  �X  B�    ��Dj                      �4  �X  B�    p	��Dj          �aG�        �4  �X  B�    ���Dj          ?��        �4  �X  B�    57���               ���>���              ;7���                ?�>B�\              `�8�f                ?   ?��              i�8�f            �\(?   ?5              )
�8�f            >#�
?   ?5              x	�8�f            ;��>���?,̼        ´    �7���               ���<���            