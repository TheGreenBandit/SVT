   ���     ra�                              }��                                      Ȗ0�           ��>B�]>B�]        B�    Ȗ0�           ?�3/>B�]>B�]        B�    rȖ0�           ?33(?�Q�?
>        B�    �Ȗ0�           =��s?�Q�?
>        B�    -Ȗ0�           >�̶�W
:?�         B�    Ȗ0�           ?L̻�W
:?�         B�    �Ȗ0�           <��ʾW
:?�         B�    �^֨^               ��(�?ٙ�        =��	  #^֨^               ��(�?ٙ�@�Q�    C�
>  
^֨^           ���;�(�?L̴@�Q�    B�(�  8^֨^           ?���k�?��@�Q�    B�(�  ^֨^           ���Ϳ���?L̴@�Q�    B�(�  �^֨^           ?333����?L̴@�Q�    A�
P  �n�~               �   ?�                �n�~           ?�  �                     2n�~           �fff4�  ���              �n�~           �fff����>���        �bff  V	n�~                    ��                �	��L                ��  �                 [
��L                ��  �              