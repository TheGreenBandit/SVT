   9�     ;�                              ��|(                              ´    ��|(          �u                ´    ��|(          ��                ´    ��|(          �0��                ´    ��|(          ?f                ´    ��|(          ?�d                ´    ��|(          @                  ´    ��|(          @}                ´    �Ȗ0�          �L�����>��P        B�    cȖ0�          �L�����=�G�        B�    qȖ0�          >.]����=�G�        B�    �Ȗ0�          >.]����>�x        B�  