   q��     u�                              /�v�n           @ff��3<�:�6��            0�v�n           @ff�Ffh@�V/��z�          C�v�n           @��?��3<�:�6��            Q�v�n           @���Ffh@�V/��z�        