   9��?                                     ��yLp               @�31>.|<#�
        