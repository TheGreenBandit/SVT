   Pѫ     ?�                              �	�0�>                                     �	�0�>               ����                  F	�0�>               �334                  �	�0�>               >���                  =
�0�>               ?L��                  �	ky^�            �\)?z�J=����F            �ky^�           >�?z�J=����F            �	�0�>               ��                    �	�c��           ��  ?L�ξ�z�              V	�c��           =��˿L�̽�Q�B�fXA���      �	�c��           ���ϿL�̽�Q�B�fX�6fj      �	<���           ��  ?��ؽ��	            