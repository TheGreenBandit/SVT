   
���      m                              �!}��                                      (Ȗ0�           ��>B�]>B�]        B�    �#Ȗ0�           ?�3/>B�]>B�]        B�    H1Ȗ0�           ?33(?�Q�?
>        B�    �Ȗ0�           =��s?�Q�?
>        B�    MȖ0�           >�̶�W
:?�         B�    :/Ȗ0�           ?L̻�W
:?�         B�    4"Ȗ0�           <��ʾW
:?�         B�    V7�v'&          @   �0(�@�  ��      ?�    &�v'&          @!G��  A�  �      ?�  