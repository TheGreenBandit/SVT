   �O�     8�                              �P���           >��?\%            �4    {P���           ��� ?\%            �4    P���           ���	?\%���        �4    	P���           >#�
?\%��=p        �4    �P���           >#��c���\         �4    )P���           >B�]>�Q���=p        õ�   �P���           �B�]�c���\(        �4    �P���           >��?z�4           �4    �
P���           ����?\%<#׀        �4    �P���           �\,�nq��p�        �4    X
P���           �\,>B�z��p�              	P���           ��z�nq��p�        �4    9P���           >�\(�np��p�        �4�  ���Dj       	                   ��  ´    q
��Dj       
                   ��  ´    ���Dj                          ��  ´    	��Dj                          ��  ´    
P���           >��np��p�        �4�  b
Ȗ0�           �(��?(��?\0        B�    �Ȗ0�           ?=p�?(��?\0        B�    ���Dj       	   �aG�2�          ��  ´    ���Dj       
   �aG�2�          ��  ´    ���Dj          �aG�2�          ��  ´    ��Dj          �aG�2�          ��  ´    �Rf�               �?��>Ǯ        �4    D�8�f                ��z�?.u    ´        ���9�                ���?h��              ���9�            <#ֺ?Y���ǭ�        �4  