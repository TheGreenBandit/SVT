   =��\                                      �}��                =�\(<��
�@            !j�&�           ��G��z�            B�    [j�&�           >.{�z�            B�    ]�k0       	    ����                B�    -�k0       
    ����                B�    b�k0           ����                B�    T�k0           ����                B�    pV���                �37>k�            