   �O�                                      ��)=�               ��G���
7              �
�)=�               >��ɿ�
7        �4    :�)=�               =�׫��
7        ´    �)=�               ���l��
7        B�    ��)=�               ���l��
7        B4    �)=�               ���l��Q���          ��)=�           >������
7        �T  