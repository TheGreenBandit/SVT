   �wb                                      q�wb                                A�    X�wb                                B     m�wb                                Bp    ��wb                                B�    W�wb                                B�  