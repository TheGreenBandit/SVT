   ,��.Q     q�                              D:�           �ff]?�>���        ´    'D:�           �ff]?��K>���        ´    �D:�           �ff]?#�>���        ´    �D:�           �ff]=#�>���        ´    �D:�           �ff]�\$>���        ´    �D:�           �z�=��3,>���    ��  ��    �D:�           �z�=��Q�>���    ��  ¯�u  �D:�           �Y���(�>���    ��  �3(�  mD:�           ��fe�"�]>��@    ��  ���  6D:�           =u�(Q�>��@    ��  7�P   �	D:�           ?\%�p�>��@    ��  B   kD:�           ?s3*� ��>�{    ��  B�G�  D:�           ?����) >��@    ��  B���  �D:�           ?���z�T>��@    ��  B���  rD:�           ?�G���G�>��@    ��  B���  �D:�           ?��>Z>��@    ��  B���  DD:�           ?p��??��>��@    ��  B���  �D:�           ?p��?���>��@    ��  B���  �D:�           ?p��?���>��@    ��  B���  jD:�           ?#�@p�>���    ��  C!  �D:�           <��0@z�>���    ��  C6!  �D:�           ��@��>���    ��  CL�.  `D:�           �z�?���?B��¦      C4!  �D:�           <��*?���?B��¦      C4!  �D:�           ?z�?���?B��¦      C4!  5D:�           ?z�?}p�?���hp�@@  C4!  D:�           <#�Z?}p�?���hp�@@  C4!  �D:�           �\$?}p�?���hp�@@  C4!  �D:�           �Q�|?8Q�?O\L?c� Brp�C���  ~D:�           �J=h>�=;?O\L�G
 ?*@C���  D:�           �O\ ����?T{�G
 ?*@C���  �D:�           �O\ �p��?T{�G
 ?*@C���  �
D:�           �ff\���?T{�G
 ?*@C���  �D:�           �O\ ��?T{�G
 ?*@C���  �D:�           ���� ��?T{�E�R?��C��  dD:�           =L���,(�?T{�E�R?��C���  	D:�           ?z��z�?T{�E�R?��Cʐ�  �	D:�           ?h������?T{�E�R?��C֐�  PD:�           ?ff^��G�?T{�E�R?��C��  {D:�           ?ff^�0��?T{�E�R?��C��  D:�           ?ff^�W
l?T{�E�R?��C��  LD:�           ?ff^>�p�?T{�E�R?��C��  �D:�           ?ff^>�p�?T{�E�R?��C��  <	D:�           ?ff^?^�>?(���E�R�{p�C��