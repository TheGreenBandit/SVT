   �%��     ��                              k�c"               >\(>�31        �6    ���X       	   �p                ´    ���X       
   �p                ´    ���X          �p                ´    ��X          �p                ´    �7���               �p�ؽu              8	Ȗ0�          �B��?�=k>�        B�    	
Ȗ0�          >�=[?�=k>�        B�    �
��X       	   ���                ´    ���X       
   �(�                ´    �	��X          ���                ´    
��X          �(�                ´    �
�8�f            =#�
?��=�G�              m�8�f           ���
�}p~?
=m              �����                                      �����           =L��?��A��         �4    �����               ?��A����        ô  