   
����     41                              �s��               �aG�                  ��B�,       	   �W
>                ´    ��B�,       
   �W
>                ´    ��B�,          �W
>                ´    ��B�,          �W
>                ´    ��B�,          ��G����ο�p�        ´    ��B�,          ��G���3.��p�        ´    ��B�,          ?��R��3.��p�        ´    ��B�,          ?��P�336��p�        ´    ���g-                @k���  �4  È  B�  