   c"��    q�                              X�            ��                        >�            ?�                        ��            =���?� ?�                ��            =���@  ?���              e�            =���@&fe?�fg              ��            =���@331?�               �            =���@?��?���              ��            =���@L��?ٙ�              ��            =���@_��?ٙ�              ��            =���@s3-?�fh              ��            =���@���@��              �
�                    @�              