   �$�     �                              zt_3�          >L���  � ��´          