   	�O�     `�                              �8��               �����Q        ´    ���Dj       	   ����                ´    ���Dj       
   ����                ´    @��Dj          ����                ´    M��Dj          ����                ´    G��9�               ����?J=���            E{��
                ����#��            L��<              @�              C4    [L��<              ��                  