   �$�                                      <�$�                                ��    _�$�                                �H    d�$�                                    A�$�                                ��    S�$�                                ��    *�$�                                �    ��$�                                �/    }�$�                                �H    z�$�                                �a    j�$�                                �z    &�$�                                É�    �$�                                Ö    N�$�                                â� 