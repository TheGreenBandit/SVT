   @�     W��                              ��3�           ?�35��fe@                 ��3�           ������fe@                 P�!�               �QG�?L��        ´    P�!�               �!G�?L��        B�    >]��                �@  @^y        C4    	��           ��`��fg?p��C4      B�    ��           @G���fg?p��C4      B�    ���                �   @W�              �M:-            ?��(�@)��C|��  A�fh  +�z            ?�34�32@  ´      B�    �i}�               �0�*?�G�        C4    �r`�               �` ?�p�        C4    /S~�               �-��?�
D              4�|F�                �2�?���        C4    ;��U            ���A�2~?���        C4    6�p��            >����2~?�        C4    H�r`�               �#��?�p�        C��   K#*�+            �334�'��?L��        C4    LP��                �+�(?���        C4    M��           ��z���G�?p��    ��C4  