   9��?    L�                              H_�d           ��@g�ӽ�\(C�� ´  �    H_�d           ���@1�G        ´  �    H_�d           ��Rl@
�=L��    ´  ��    	H_�d           >v?�����\(    ´  A�    H_�d           �ǭ�@a�D��    ´  �    �H_�d           ����@O����\(    ´  �4    �H_�d           ��@+�὏\(    ´  �F    :H_�d           ��
,@�὏\(    ´  C    H_�d           �W
"@�
��\(    ´  C�    xH_�d           �u�t@s2w��\(    ´  C�    H_�d           �u�t@s2w��G��6\)�  C�    H_�d           �u�t@O�F���5 �4  C�    �H_�d           �u�t@o���4 �4  C�    H_�d           �u�t@o�>�<�4     C4    H_�d           �u�t@O�F>�p��5 ô  C�    PH_�d           �u�t@l(:>�z��6Q���  C�  