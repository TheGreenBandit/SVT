   ��     P�M                              �
Qp��                    ?�                
Qp��            >���    ?�                BQp��            �      ?�                �
Qp��            �ffh    ?332              �
Qp��            ?ffg    ?332              AQp��            ?ffg    >���              {
Qp��            �ffh    >���              1Qp��            ����    ?�34              �
Qp��            >���    ?�34              �
Qp��            ��      ?ٙ�              v
Qp��            ��  @��@l���   �   ®    <Qp��            ��  @��@,��´  ��  ®    Qp��            ��  @��@l��´  ��  ®  