   ͓��     �w                              ept�               >�G�            @@    f:��E               ��>���              g���                   >�
9�#�
        