   v*�                                     �v*�                           �        �v*�                           B      