   �]�     �G�                              �.�]�                            ��        �@ȟ�                                      ��]�                            �         ;@�]�                            �p        �E�]�                                     �B�]�                            A�        ->�]�                            B         �=�]�                            Bp        �2�]�                            B�        ��8�f                �
=p>��               #A�8�f               �
=p=u�@              �F�8�f           ��  @��L�A�            oF�V                �`?��    ô        �E7���           ?����?��    ��33      d?7���           ��\���?5¤    ��33      �E7���           ���P���$>W
�    ��33      +7���           ?���������j    ��33      YC�M:-           ��\(>\*=�Q�B�  ¥���)4  K.�M:-           ?�=p>\*=�Q�B�  £��;?�  F�V            �J=i�`?��    ô        /D�V            ?&fa�`?��    ô        �1�V            ?&fa�`>���    ô        55�M:-           ��[�>#�
?� 
C1  �4��~h�