   �O�                                     x��               @_��?�f_              ��M:-           ����?�  @     A�
BB
z�  ��M:-           ����?�  ?���  A�
BB
z�  ��M:-           ����?�  =�̣  A�
BB
z�