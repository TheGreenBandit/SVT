   2,��     ��;                              �	���                <#�
��Q�              6%Z_�       	   �aG�                ´    �%Z_�       
   �aG�                ´    �%Z_�          �Z                ´    �	%Z_�          �Z                ´    �	���v           =��aG�>k�!´            ����v           >���aG�>k�!´            >	���v           ?��ϾaG�>k�!´            ����v           ?����aG�>k�!´            �	���v           ?�������L��´            �	���v           ?�p�����B�]´            �	���v           =�����B�]´            E	���v           =�����#�
´            �	���^              @@              C4    ����^              �   @5�A`      C4  