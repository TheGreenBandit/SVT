    ���     &�                              ���Dj       	                       B�    R��Dj       	   >�=q                B�    !��Dj       	   ��=r                C�    z��Dj          ��=r                C�    s��Dj          �
=l                C�    c��Dj          3�                  C�    ���Dj          >�=t                C�    4��Dj          ?�                B�    xȖ0�           ���?�  ���<#�
    B�    �Ȗ0�           ?�?�  ���<#�
    B�    ~��E�                �Qhh>m�~�   Ç        07���                >�y>� A�            ��8�f                ��Q�>Ǯ��             �8�f                �!G�>�(�A          