   c"��                                     �            ��                        �            ?�                        �            =���?� ?�                4�            =���@  ?���              #�            =���@&fe?�fg              P�            =���@331?�               Z�            =���@?��?���              ��            =���@L��?ٙ�              [�            =���@_��?ٙ�              v�            =���@s3-?�fh              ��            =���@���@��            