   9��?     �                              � �3�           B�u��陜�=�               �3�           A�39=z��(�          