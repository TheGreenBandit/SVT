   �O�                                      cGY^&                �ٙ�����              VGY^&                ?�  ����              b%Z_�       	    @~                ´    f%Z_�       
    @~                ´    j%Z_�           @~                ´    o%Z_�           @~                ´  