   �D�                                      *
<
�           �!G�<�� ����¶36B�  �     �<
�           �!G�<�>¶36B�  �     �<
�           �!G�<�>�{¶36B�  �     )<
�           �!G�<�>�f�¶36B�  �     <
�           �!G�<�?��¶36B�  �     I<
�           ?�<�?��¶36B�  �4    �<
�           ?�<�>�G�¶36B�  �4    �<
�           ?�<�>�=�¶36B�  �4    
<
�           ?��=�Q�=�Hf¶36B�  �4    �
<
�           ?�X<��#�:¶36B�  �4    f<
�           54  ?u >Ǯ>��    �4    �<
�           54  ?Y��>�¶��    �4    �<
�           �#�:?=p�?)��    �4    �<
�           <�������>�f�Å��    �4    <
�           <�������>���Å��    �4    �<
�           <�������>\�Å��    �4  