   �Z�     @�                              `}��               =�\*=����)          �Ȗ0�           ?�  >��>�\@        B�    �Ȗ0�           ��=p>�넽L�        B�    �Ȗ0�           ?��>�넽L�        B�    	Ȗ0�           ���Q>��>�\@        B�    w��                ?�Q�=��4            w��                >�=��4            w��                ����=�G��4            �w��            ?(��?���=R��  @�        �w��            �(��?���=�q��  ��        ���Dj       
   ��=q                ´    ���Dj          ��=q                ´    ���Dj          ��=q                ´    ���Dj       	   ��=q                ´    n�v'&              �P��@�f`��            ��v'&              �'
A�\K�,          