   
���    ���                              E6}��                                     6Ȗ0�         ��>B�]>B�]        B�    �4Ȗ0�         ?�3/>B�]>B�]        B�    �6Ȗ0�         ?33(?�Q�?
>        B�    R6Ȗ0�         =��s?�Q�?
>        B�    �5Ȗ0�         >�̶�W
:?�         B�    �7Ȗ0�         ?L̻�W
:?�         B�    C6Ȗ0�         <��ʾW
:?�         B�    Q5�v'&                      ��      ?�    H7�v'&              �p  A   �      ?�  