   .���     a�                              /�y�e           ���U�3���
#              ��y�e           ���U�3�>��h              7�y�e           ���U��
�>��h              &�y�e           ���U@%�>B��              8�y�e           �#���3�>���    <��
      �y�e           ?����3�>���    <��
      C�y�e           ?����&f�>���    <��
      �y�e           ?���@3.>���    <��
    