   ��    <�                              �Qp��                    ?�                *Qp��            >���    ?�                iQp��            �      ?�                <Qp��            �ffh    ?332              EQp��            ?ffg    ?332              +Qp��            ?ffg    >���              )Qp��            �ffh    >���              Qp��            ����    ?�34              0Qp��            >���    ?�34              HQp��            ��      ?ٙ�              �Qp��            ��  @��@l���   �   ®    -Qp��            ��  @��@,��´  ��  ®    Qp��            ��  @��@l��´  ��  ®  