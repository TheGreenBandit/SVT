   �O�                                     v�3�               �������              [�y�e               ���A��z�              ��y�e               ���A�#�              r�y�e               ���A>\'            