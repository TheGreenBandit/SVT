   �%��    p��                              "���               >�G��\%              6O|y�                ?
~�>ܬ              7��               >���>���              8s���               ��\@��        �2    9[�3           �&fa>��>�(�              :g��           ?�>�fa>�G�        �4  