   	ց                                      ����v            �
9?�p�>�K�´            ����v            �?��?˅">���´            =���v            ?@ 0?Ǯ?*�´            k���v            ?
9?�p�>�K�´            �1A�           �
=m?�p�?aG�        B�    �1A�           ?�?�p�?aG�        B�    �1A�           ?��>#�7?z�        B�    }1A�           ���>#�7?z�        B�    j}��                   ?
=m            