   c"��   �>�                              �*(�E�                @�
?xQ�C4            !(�E�            �   �\*?xQ�C4      �4    [,(�E�            @@  ?�X?xQ�C4      ³��  \*(�E�            ����@�Q�?xQ�C4      B� )  /"���^          ?
=m@�fc�\(    ��  �4  