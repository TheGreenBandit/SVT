   {~V�                                      3{~V�                               �4  