   c"��                                      �	�oX/           ?�  A   �334              )
�oX/           ?�  A�  �334              p
�oX/           ?�  A�  �334              �
�oX/           ?�  B  �334            