   KlV�                                      �7���            2�      ?�fh              �7���            ����L��>L���f�          N7���            2�  ?   ?�fh              :7���           ����?   ?�fh              37���           >���?   ?�fh              V7���            ?���L��>L���f�        