   q��     �                              W}��                   =�Q�ff]          YȖ0�            ���W?!G�=��%        B�    ZȖ0�            ?��?!G�=��%        B�    [Ȗ0�            >X?�=e>��h        B�    \Ȗ0�            ���?�=e>��h        B�  