   �O�     &�                              r��L                ?��>�f`        ´    H��L                ����>�f`        ´    G	��L                �n�>�f`        ´    �	��L                �n�>�fa´  ��  ´    ~	��L                �W
J>�fa´  ��  ´    E	��L                ?(�>�fa´  ��  ´    ���L            2�  ?(��>�fa´  ��  Ç    	��L            2�  �B�f>�fa´  ��  Ç    d	��L            2�  �5>�fa´  ��  Ç    =	��L            2�  �p��>�fa�4  ´  Ç    �	��L                ?330>�f`�4  Ç  Ç    �	��;#       	   ��                ´    �	��;#       
   ��                ´    w	��;#          ��                ´    �	��;#          ��                ´  