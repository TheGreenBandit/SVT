   ��\�                                      �.�                =�Q�=���              ���Dj       	   �u                ´    ���Dj       
   �u                ´    ���Dj                              ´    b��Dj          ?��                ´    ���Dj          ?��                ´    ���Dj          �
9                ´    ���Dj          �
9                ´    �O{Q�           ����?�G�>���B,      C4    �O{Q�           ����@�>��B,      C4    �O{Q�           �W
m@�	��ՠB,      C4    2�5�V            �ff]�}p��L��        B�    ��5�V            �ff]�}p��z�        B�    \�5�V            ?ff]�}p��z�        B�    ��5�V            ?ff]�}p��^�I        B�    FO{Q�           >L̠@�	��ՠB,      C4    7O{Q�           >�=[@�>��B,      C4    �O{Q�           >�=[?��
>�z�B,      C4  