   C*�f                                      3�܇                                     C�܇                                     E�܇       
                              D�܇       	                            