   �q�4     c�                              �7l�               ��Q���              ��܇       	   ����                      ��܇       
   ����                      ��܇          ����                      ��܇          ����                      ��%�;            =u@��?0��    ´        ��%�;            =u@��O�u�\A�  ´        ��%�;            ��\ @I�>?  
�#�
´  B�    ��%�;            ��\ ?L�v?  
�#�
´  B�    ��%�;            ��\ ���z?  
�#�
´  B�    ��%�;            ��\ �� (?  
�#�
´  B�    ��%�;            �S��f�?  
�#�
´  B�    ��%�;            ��3)��ܽ��`�#�
�4 B�    ��%�;            ��3)?�|���_�#�
�4 B�    ��%�;            ��3)@�[�>���#�
�4 B�    ��%�;            ?�fv@I�>?  
�#�
´  ´    ��%�;            ?�fv?L�j?  
�#�
´  ´    �%�;            ?�fv�� �?  
�#�
´  ´    �%�;            ?�fv�s3�?  
�#�
´  ´    �%�;            ?�fv��f�?  
�#�
´  ´    ��%�;            >B���ٙr>�\D�#�
B�  �13.  ��%�;            ?� @�Go���_�#�
�4 ´    �%�;            ?� ��h���`�#�
�4 ´    ��%�;            ?� @�z����`�#�
�4 ´    ��%�;            ?� ��gN���`�#�
�4 ´    ��%�;            >B���ٙr?� �#�
B�  �13.  ���^              A1�|����        �4    ����^              @�[�?���Au�v    �4  