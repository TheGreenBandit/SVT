   �)��    ��=                              *�           ����    �B�\        �4  