   �O�    NĮ                              �t�-�               >�=r�B�U        C4  