   ����                                      n�            �����334?���A�f�          �n�            >��̿334?���A�f�          <wMl]           �����33?334?�fi          0wMl]           ����33?334?�fi          QwMl]           ?�35�33?334?�fi          �JF��            �9���,��?ffh��  A�  ´ff  �wMl]           ����@l��@331@���          �wMl]           ����@�3*@���Aff          �wMl]           ?��@�3#@���A� ��fi�/L�  \wMl]           >���A.fi@  A\�޿�fi�/L�  �wMl]           >L��AQ��?336A�ο�fi�/L�  �wMl]           >���Ax ����A�ο�fi�/L�