   �O�     	��                              ���g-               �#�                  ���g-               ?0��                  ��Dj       	   �:�A                ´    0��Dj       
   �:�A                ´    3��Dj          �:�A                ´    :��Dj          �:�A                ´  