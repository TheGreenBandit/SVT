   �O�     \CA                              ����k                �L��?!G�        B�    ���Dj       	   �Q�        �4      B�    @��Dj       	   ��38                B�    R��Dj       	   ���                B�    ��Dj       
   ��                B�    z��Dj       
   �G�                ´    ���Dj       
   ����                B�    ���Dj          ����                B�    ���Dj          ���B                C�    :��Dj          ���
                C�    ���Dj          ��Q�                B�    7���                ��\&�#�:              �
�8�f                �� >p              !?�                                      �8�f               ?�3+?z�              ��8�f               ��Q�?z�            