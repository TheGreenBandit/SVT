   c"��                                     �	�i�               �C3>?ffh              �	�,�           @�  �@                    �	�,�           ��  �@                  