   �Z�     R��                              +}��               =�G�>8Q�@]p~          �
Ȗ0�           ?�  >��>�\@        B�    �
Ȗ0�           ��=p>�넽L�        B�    �
Ȗ0�           ?��>�넽L�        B�    �
Ȗ0�           ���Q>��>�\@        B�    R
��Dj       
   ����                ´    �
��Dj          ��=q                ´    Z	��Dj          ��=q                ´    
��Dj       	   ��G�                ´    $=f�M           �xQ�>�Q�>�fb  ´        �
�E	               ?ٙ���֢´            ��E	           >�\)?ٙ���֢´            W
�E	           ���?ٙ���֢´            �
�E	           ���?ٙ�>8Q�´            �E	           ��  ?ٙ�>8Q�´            U�E	           >��?ٙ�>8Q�´            �
7���           �#�����\)              ��y�e                ��`<���B�          