   �]�                                      D�]�                           ��        dȟ�                                     E�]�                           �         G�]�                           �p        _�]�                                    ��]�                           A�        n�]�                           B         [�]�                           Bp        ��]�                           B�        ^�8�f               �
=p>��               k�8�f               �
=p=u�B              ��8�f           ��  @��L�A�          