   �]�                                      ��]�                                �p    ��]�                                ��    �	�]�                                �4    y	�]�                                �p    	�]�                                    "�]�                                ´    ��]�                                ��    *	�]�                                ��    �	�]�                                �    �	�]�                                �    }	�]�                                �     �	�]�                                �/    	�]�                                �>    9�]�                                �M    =	�]�                                �\    m	�]�                                �k    �	�]�                                �z    ��]�                                Ä�   
�]�                                Ì    �	�]�                                Ó�   ��]�                                Û    �	�]�                                â�   �	�]�                                ê    B�]�                                ñ�   U	�]�                                ù  