   ��.Q   ,�                              �	]
��           ��\(?���� <�          �����           =u�j�E�33-        B�    �%&�N           >L���   �O\!        B�    �	�)�=           ?   �@  �L��        B�    �	�D�            ?��@(�>���k�!<#�@���  �	�D�           ?
=m�L��>�            