   �l     M�                              ���Dj       	                   A`  B�    ���Dj                          A`  B�    ���Dj          >�             A`  B�    ���Dj          >�            A`  B�    ���Dj          ?=p�            A`  B�    7��Dj          ?��            A`  B�    ���Dj          ��             A`  B�    ���Dj          ��            A`  B�    ���Dj          �:�A            A`  B�    ���Dj          �z�>            A`  ´    ���Dj       	   �k�             A`  C�    ���Dj       	   >aG�            A`  B�    ��8�f                ?(�?��              ��8�f                ?.z>�G�              ��8�f                ??��>�\,              ��8�f                >�3<>��DB0            ��8�f                =���>��TA�            ��8�f                ��H>��T�.�          �7���            �#�
=#�
��G�A�            ��8�f           ��fd<�ت<�·�.�          ��8�f           ?�fk5P  <�·�.�          ��8�f       	    ?
=u��Ӣ=L�X�.�          ��8�f       	    �\<��r=L�X�.�        