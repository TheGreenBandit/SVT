   B��     %
?                              �� �^                ��  �#�
              5D:�            �G����?L����  C�  C�    �=f�M            �\'��|?.��P  B�        �Ȗ0�           �W
>����B�]        B�    �Ȗ0�           >L�Ϳ���B�]        B�    s�8�f                @�ž\(              ��8�f                �8��>��T��            �%Z_�       	   ��G�                B�    �%Z_�       
   ��G�                B�    �%Z_�           ���                B�    �}��                ��>���              �D:�            �G��z�?L����  C� C�    ,D:�            ?G��z�?L��CK  C���C�    YD:�            ?G��}p�?L��CK  D�C�    �=f�M            >���|?.��P  B�        %Z_�           ���                B�  