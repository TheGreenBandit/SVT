   ���     �                              z}��                                      �Ȗ0�           ��>B�]>B�]        B�    Ȗ0�           ?�3/>B�]>B�]        B�    �Ȗ0�           ?33(?�Q�?
>        B�    �Ȗ0�           =��s?�Q�?
>        B�    �Ȗ0�           >�̶�W
:?�         B�    �Ȗ0�           ?L̻�W
:?�         B�    �Ȗ0�           <��ʾW
:?�         B�    ��v'&           @�  �0(�@�  ��      ?�    ��v'&           @���  A�  �      ?�    D*�v'&           @���`  Bp��      ?�  