   �                                      �D:�           �Q눿0��?�
<        ´    �D:�           �Q눿�?�
<        ´    �D:�           �Q눿��?�
<        ´    �D:�           �Q���?�
<        ´    �D:�           �  ��B?�
<              �D:�           =L���B?�
<              �D:�           ?�N��B?�
<              �D:�           ?L̺�z�?�
<        B�    �D:�           ?L̺�˅?�
<        B�    �D:�           ?L̺��\(?�
<        B�    �D:�           ?L̺�+�$?�
<        B�    �D:�           >���3H?�
<        C4    �D:�           <�ժ��3H?�
<        C4    �D:�           ����3H?�
<        C4    �Ȗ0�           ��R @z�?L��        B�    �Ȗ0�           >�\@z�?L��        B�  