   �"�                                     ,ky^�           �   2�  2�                B(ky^�           �   2�  2�                �(ky^�       
    �   2�  2�                }+ky^�       	    �   2�  2�              