   �l                                      }��Dj       	                   A`  B�    ���Dj                          A`  B�    ��Dj          >�             A`  B�    ���Dj          >�            A`  B�    :��Dj          ?=p�            A`  B�    ���Dj          ?��            A`  B�    ���Dj          ��             A`  B�    �
��Dj          ��            A`  B�    ���Dj          �:�A            A`  B�    ���Dj          �z�>            A`  B�    ���Dj       	   �k�             A`  B�    ���Dj       	   >aG�            A`  B�    ��8�f                ?(�?��              ~�8�f                ?.z>�G�              c�8�f                ??��>�\-              ��8�f                >��>ǮA�            ��8�f                ����>uA�            �8�f                ��H>��T�.�        