   @�     �:[                              �!               ��p�?z�        B�  %B�<           >�(�    @           C��   ��!               ��p�@6fd        B�  a�!               ��p�@tz�        B�  8�^�R           ��  �330@���        B�    r�!               ��?z�        B�  E#�!               ��@6fd        B�  ��!               ��@tz�        B�