   ��                                      ����                ?�fh    A���          ����            �� �0��?z�GA*fn    C3    ����            >���0��?z�GA*fn    C3    ����            >���0��?��
A*fn    C3    ����            �� �0��?��
A*fn    C3    ����            �� �0��?�=qA*fn    C3    ����            >���0��?�=qA*fn    C3    ����                ��fg>���A���        