   �D�                                      ��D�           ?�                       ��D�               �L��                  b�D�           ?� �L��                  �JF��               �L��?332        ´    �JF��           ?� �L��?332        ´    �JF��           ���˾���>L��B�      ´    �JF��           ���˾���?@  B�      ´    JF��           ?�(辙��?J=p´      ´    tJF��           ?�(辙��?J=p´      ´    �JF��           ?�(辙��>k�>´      ´    �D:�           �W
@?�V?B�^�Qk2�  �3��  �D:�           >�=q?�V?B�^�Qk2�  �3��  �D:�           ??��?�V?B�^�Qk2�  �3��  �D:�           ?���?�V?B�^�Qk2�  �3��  �D:�           ?�
5�z�?B�^����4   7�    �D:�           ?Tz��z�?B�^����4   7�    �D:�           >k�&�z�?B�^����4   7�    zD:�           ��p��z�?B�^����4   7�  