   c"��     G�                              �|{B           A`      �Y        Cx    �|{B           A`  >8Q�A���        C�    �|{B           A`  >�=qBz�        C��   �|{B           A`  >�p�BJ�        C�    �|{B           A`  >�G�B�B�        C�    �|{B           A`  >�B�B�        C��   �|{B           A`  ?\%B�B�        C�    �����           A]�?u�|B�]        �L  