   ���     </�                              _��M                                A�    t��M                                A�    ��M                                B4    ��M                                Bh    ���M                                B�    ���M                                B�    ���M                                B�    ���M                                B�    ���M                                C    ��M                                C    ���M                                C    ���M                                C+    8��M                                C8    ���M                                CE    ���M                                CR    ���M                                C`    ���M                                Co    ��M                                C~    ���M                                C�    ���M                                C�    
��M                                C�    ��M                                C�    ���M                                C��   ���M                                C��   	��M                                C�� 