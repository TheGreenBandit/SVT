   2,��     "�X                              E���                <#�
��Q�              G%Z_�       	   �aG�                ´    ;%Z_�       
   �aG�                ´    1%Z_�          �Z                ´    "%Z_�          �Z                ´    J���v           =��aG�>k�!´            K���v           >���aG�>k�!´             ���v           ?��ϾaG�>k�!´            P���v           ?����aG�>k�!´            N���v           ?�������L��´            ���v           ?�p�����B�]´            M���v           =�����B�]´            H���v           =�����#�
´            ��v'&          =�������@���C          