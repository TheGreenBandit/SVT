   ���     H<�                              �}��                                      C	Ȗ0�           ��>B�]>B�]        B�    �	Ȗ0�           ?�3/>B�]>B�]        B�    �	Ȗ0�           ?33(?�Q�?
>        B�    
Ȗ0�           =��s?�Q�?
>        B�  