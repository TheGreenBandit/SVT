   	��     ]�^                              �
��            >\(��  ���	        B�    �
Md�            ��������?�=oB��    ��    �
Md�            >L�̾���?�=oB��    ��    �
�V            >���?   =L���ff          �
�V            ��=r?Y��2   @�34    �3    �k0       
   �#�
                C�V  �k0       	   �#�
                C�V  F	�k0          �#�
                C�V  �
�k0          �#�
                C�V